* NGSPICE file created from tt_um_urish_charge_pump.ext - technology: sky130A

.subckt tt_um_urish_charge_pump clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VAPWR VGND VDPWR
X0 vout.t3 w_20072_2496.t2 w_20072_2496.t3 vout.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=40
D0 stage3.t1 vout.t0 sky130_fd_pr__diode_pd2nw_11v0 pj=4e+06 area=1e+12
X1 ua[0].t3 VGND.t3 VGND.t4 ua[0].t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=40
D1 stage1.t1 stage2.t0 sky130_fd_pr__diode_pd2nw_11v0 pj=4e+06 area=1e+12
X2 clka clk.t0 VGND.t1 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 clkb.t1 clka VGND.t2 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
D2 VAPWR.t3 stage1.t0 sky130_fd_pr__diode_pd2nw_11v0 pj=4e+06 area=1e+12
X4 VGND.t5 vout.t1 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X5 ua[0].t1 ua[0].t0 w_20072_2496.t1 w_20072_2496.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=40
X6 stage1.t2 clka.t0 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X7 VAPWR.t1 clk.t1 clka VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
D3 stage2.t1 stage3.t0 sky130_fd_pr__diode_pd2nw_11v0 pj=4e+06 area=1e+12
X8 stage2.t2 clkb.t0 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X9 VAPWR.t2 clka clkb.t2 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X10 stage3.t2 clka.t1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
R0 w_20072_2496.t2 w_20072_2496.t0 644.312
R1 w_20072_2496.t1 w_20072_2496.t2 660.668
R2 w_20072_2496.t2 w_20072_2496.t3 660.264
R3 vout.n21 vout.n15 8605.04
R4 vout.n18 vout.n16 8605.04
R5 vout.n19 vout.n15 3489.23
R6 vout.n20 vout.n16 3489.23
R7 vout.n22 vout.n14 1652.71
R8 vout.n17 vout.n14 1652.71
R9 vout.n17 vout.n13 1652.71
R10 vout.n23 vout.n22 1451
R11 vout.n5 vout.n2 741
R12 vout.n9 vout.n2 741
R13 vout.n9 vout.n3 741
R14 vout.n24 vout.t3 660.414
R15 vout.n8 vout.t0 323.575
R16 vout.n6 vout.n5 236.839
R17 vout.n23 vout.n13 167.992
R18 vout.n8 vout.n7 151.427
R19 vout.n4 vout.n0 146.447
R20 vout.n4 vout.n1 146.447
R21 vout.n10 vout.n1 125.314
R22 vout.n11 vout.n0 123.569
R23 vout.n5 vout.n4 46.2505
R24 vout.n10 vout.n9 46.2505
R25 vout.n9 vout.n8 46.2505
R26 vout.n3 vout.n1 46.2505
R27 vout.n2 vout.n0 46.2505
R28 vout.t0 vout.n2 46.2505
R29 vout.n15 vout.n14 37.0005
R30 vout.n16 vout.n13 37.0005
R31 vout.n6 vout.n3 29.6199
R32 vout.t0 vout.n6 14.7834
R33 vout vout.n24 8.20169
R34 vout.n12 vout.n11 2.16948
R35 vout.n24 vout.n23 1.75703
R36 vout.n11 vout.n10 1.74595
R37 vout.n22 vout.n21 1.54217
R38 vout.n18 vout.n17 1.54217
R39 vout vout.n12 1.09447
R40 vout.n21 vout.n20 0.917376
R41 vout.n19 vout.n18 0.917376
R42 vout.n20 vout.t2 0.626126
R43 vout.t2 vout.n19 0.626126
R44 vout.n12 vout.t1 0.404364
R45 stage3.n9 stage3.n2 741
R46 stage3.n6 stage3.n2 741
R47 stage3.n7 stage3.n6 741
R48 stage3.n5 stage3.t0 323.575
R49 stage3.n9 stage3.n8 236.839
R50 stage3.n5 stage3.n4 151.427
R51 stage3.n3 stage3.n0 146.447
R52 stage3.n3 stage3.n1 146.447
R53 stage3.n10 stage3.n1 142.268
R54 stage3.n11 stage3.n0 135.774
R55 stage3 stage3.t1 68.9393
R56 stage3.n10 stage3.n9 46.2505
R57 stage3.n6 stage3.n3 46.2505
R58 stage3.n6 stage3.n5 46.2505
R59 stage3.n7 stage3.n1 46.2505
R60 stage3.n2 stage3.n0 46.2505
R61 stage3.t0 stage3.n2 46.2505
R62 stage3.n8 stage3.n7 29.6199
R63 stage3.n8 stage3.t0 14.7834
R64 stage3.n11 stage3.n10 4.8005
R65 stage3.n12 stage3.n11 4.61856
R66 stage3.n12 stage3.t2 2.68428
R67 stage3.n13 stage3.n12 1.52064
R68 stage3 stage3.n13 0.1255
R69 stage3.n13 stage3 0.063
R70 VGND.n29 VGND.n22 2.10485e+06
R71 VGND.n60 VGND.n41 2.0614e+06
R72 VGND.n41 VGND.n30 1.98293e+06
R73 VGND.n30 VGND.n29 338800
R74 VGND.n75 VGND.n22 184568
R75 VGND.n23 VGND.n12 50298.8
R76 VGND.n32 VGND.n30 18002.7
R77 VGND.n30 VGND.n25 18002.7
R78 VGND.n60 VGND.n26 17143.9
R79 VGND.n60 VGND.n43 17143.9
R80 VGND.n41 VGND.n40 13280.2
R81 VGND.n44 VGND.n42 9131.66
R82 VGND.n56 VGND.n42 9131.66
R83 VGND.n31 VGND.n22 9057.83
R84 VGND.n76 VGND.n75 8496.85
R85 VGND.n54 VGND.n53 7810.05
R86 VGND.n75 VGND.n74 2792.53
R87 VGND.n73 VGND.n25 2624.6
R88 VGND.n69 VGND.n25 2624.6
R89 VGND.n69 VGND.n26 2624.6
R90 VGND.n73 VGND.n26 2624.6
R91 VGND.n62 VGND.n43 2624.6
R92 VGND.n62 VGND.n44 2624.6
R93 VGND.n66 VGND.n43 2624.6
R94 VGND.n66 VGND.n44 2624.6
R95 VGND.n35 VGND.n31 2624.6
R96 VGND.n35 VGND.n32 2624.6
R97 VGND.n39 VGND.n31 2624.6
R98 VGND.n39 VGND.n32 2624.6
R99 VGND.n56 VGND.n49 2624.6
R100 VGND.n56 VGND.n55 2624.6
R101 VGND.n51 VGND.n49 2624.6
R102 VGND.n55 VGND.n51 2624.6
R103 VGND.n78 VGND.n10 1570.81
R104 VGND.n78 VGND.n11 1570.81
R105 VGND.n79 VGND.n11 1570.81
R106 VGND.n79 VGND.n10 1570.81
R107 VGND.n21 VGND.n13 1570.81
R108 VGND.n21 VGND.n14 1570.81
R109 VGND.n17 VGND.n14 1570.81
R110 VGND.n17 VGND.n13 1570.81
R111 VGND.n68 VGND.n67 1318.44
R112 VGND.n61 VGND.n60 1219.27
R113 VGND.n60 VGND.n23 1084.89
R114 VGND.n61 VGND.n42 740.399
R115 VGND.n52 VGND.n42 740.399
R116 VGND.n104 VGND.t4 660.787
R117 VGND.t0 VGND.n12 461.221
R118 VGND.t0 VGND.n76 461.221
R119 VGND.n67 VGND.n42 400.31
R120 VGND.n54 VGND.n42 400.31
R121 VGND.n72 VGND.n27 304.565
R122 VGND.n72 VGND.n71 304.565
R123 VGND.n64 VGND.n63 304.565
R124 VGND.n63 VGND.n45 304.565
R125 VGND.n37 VGND.n36 304.565
R126 VGND.n36 VGND.n34 304.565
R127 VGND.n50 VGND.n48 304.565
R128 VGND.n50 VGND.n47 304.565
R129 VGND.n75 VGND.n23 263.846
R130 VGND.n57 VGND.n48 221.901
R131 VGND.n58 VGND.n47 220.668
R132 VGND.n71 VGND.n70 190.976
R133 VGND.n28 VGND.n27 190.381
R134 VGND.n77 VGND.n9 184.095
R135 VGND.n77 VGND.n8 184.095
R136 VGND.n80 VGND.n9 184.095
R137 VGND.n20 VGND.n19 184.095
R138 VGND.n19 VGND.n18 184.095
R139 VGND.n18 VGND.n16 184.095
R140 VGND.n53 VGND.n52 183.243
R141 VGND.n38 VGND.n37 182.732
R142 VGND.n34 VGND.n33 181.916
R143 VGND.n65 VGND.n45 180.809
R144 VGND.n65 VGND.n64 180.809
R145 VGND.n16 VGND.n15 175.812
R146 VGND.n40 VGND.n22 155.025
R147 VGND.n16 VGND.n13 146.25
R148 VGND.t0 VGND.n13 146.25
R149 VGND.n19 VGND.n14 146.25
R150 VGND.t0 VGND.n14 146.25
R151 VGND.n80 VGND.n79 146.25
R152 VGND.n79 VGND.t0 146.25
R153 VGND.n78 VGND.n77 146.25
R154 VGND.t0 VGND.n78 146.25
R155 VGND.n81 VGND.n80 129.13
R156 VGND.n18 VGND.n17 97.5005
R157 VGND.n17 VGND.n12 97.5005
R158 VGND.n21 VGND.n20 97.5005
R159 VGND.n76 VGND.n21 97.5005
R160 VGND.n10 VGND.n9 97.5005
R161 VGND.n12 VGND.n10 97.5005
R162 VGND.n11 VGND.n8 97.5005
R163 VGND.n76 VGND.n11 97.5005
R164 VGND.n82 VGND.t1 83.2145
R165 VGND.n7 VGND.t2 83.1263
R166 VGND.n29 VGND.n24 68.6903
R167 VGND.n73 VGND.n72 58.5005
R168 VGND.n74 VGND.n73 58.5005
R169 VGND.n64 VGND.n44 58.5005
R170 VGND.n63 VGND.n62 58.5005
R171 VGND.n62 VGND.n61 58.5005
R172 VGND.n45 VGND.n43 58.5005
R173 VGND.n71 VGND.n26 58.5005
R174 VGND.n27 VGND.n25 58.5005
R175 VGND.n37 VGND.n32 58.5005
R176 VGND.n36 VGND.n35 58.5005
R177 VGND.n35 VGND.n24 58.5005
R178 VGND.n34 VGND.n31 58.5005
R179 VGND.n39 VGND.n38 58.5005
R180 VGND.n40 VGND.n39 58.5005
R181 VGND.n66 VGND.n65 58.5005
R182 VGND.n67 VGND.n66 58.5005
R183 VGND.n70 VGND.n69 58.5005
R184 VGND.n69 VGND.n68 58.5005
R185 VGND.n55 VGND.n48 58.5005
R186 VGND.n55 VGND.n54 58.5005
R187 VGND.n51 VGND.n50 58.5005
R188 VGND.n53 VGND.n51 58.5005
R189 VGND.n49 VGND.n47 58.5005
R190 VGND.n52 VGND.n49 58.5005
R191 VGND.n57 VGND.n56 58.5005
R192 VGND.n81 VGND.n8 54.9652
R193 VGND.n68 VGND.n41 26.0865
R194 VGND.n105 VGND.n104 26.0302
R195 VGND.n82 VGND.n81 9.3005
R196 VGND.n15 VGND.n7 9.3005
R197 VGND.n20 VGND.n15 8.28285
R198 VGND.n104 VGND.t3 7.28674
R199 VGND.n59 VGND.n58 6.12686
R200 VGND.n83 VGND.n7 5.60682
R201 VGND.n83 VGND.n82 5.47406
R202 VGND.n74 VGND.n24 5.13619
R203 VGND.n102 VGND 4.20543
R204 VGND.n106 VGND.n105 3.8545
R205 VGND.n102 VGND.n101 2.62623
R206 VGND.n84 VGND.n83 2.49486
R207 VGND.n46 VGND.n6 1.32214
R208 VGND.n59 VGND.n46 1.27232
R209 VGND.n65 VGND.n59 1.1078
R210 VGND.n46 VGND.n28 1.1078
R211 VGND.n33 VGND.n6 1.1078
R212 VGND.n38 VGND.n33 0.817521
R213 VGND.n70 VGND.n28 0.595849
R214 VGND.n85 VGND.n84 0.56121
R215 VGND.n84 VGND.n6 0.54288
R216 VGND VGND.n106 0.365382
R217 VGND.n0 uio_oe[7] 0.32762
R218 VGND.n58 VGND.n57 0.27284
R219 VGND.n101 uio_oe[0] 0.213567
R220 VGND.n85 uo_out[0] 0.1979
R221 VGND.n86 uo_out[1] 0.1979
R222 VGND.n87 uo_out[2] 0.1979
R223 VGND.n88 uo_out[3] 0.1979
R224 VGND.n89 uo_out[4] 0.1979
R225 VGND.n90 uo_out[5] 0.1979
R226 VGND.n91 uo_out[6] 0.1979
R227 VGND.n92 uo_out[7] 0.1979
R228 VGND.n93 uio_out[0] 0.1979
R229 VGND.n94 uio_out[1] 0.1979
R230 VGND.n95 uio_out[2] 0.1979
R231 VGND.n96 uio_out[3] 0.1979
R232 VGND.n97 uio_out[4] 0.1979
R233 VGND.n98 uio_out[5] 0.1979
R234 VGND.n99 uio_out[6] 0.1979
R235 VGND.n100 uio_out[7] 0.1979
R236 VGND.n5 uio_oe[1] 0.1979
R237 VGND.n4 uio_oe[2] 0.1979
R238 VGND.n3 uio_oe[3] 0.1979
R239 VGND.n2 uio_oe[4] 0.1979
R240 VGND.n1 uio_oe[5] 0.1979
R241 VGND.n0 uio_oe[6] 0.1979
R242 VGND.n5 VGND.n4 0.13022
R243 VGND.n4 VGND.n3 0.13022
R244 VGND.n3 VGND.n2 0.13022
R245 VGND.n2 VGND.n1 0.13022
R246 VGND.n1 VGND.n0 0.13022
R247 VGND.n86 VGND.n85 0.13022
R248 VGND.n87 VGND.n86 0.13022
R249 VGND.n88 VGND.n87 0.13022
R250 VGND.n89 VGND.n88 0.13022
R251 VGND.n90 VGND.n89 0.13022
R252 VGND.n91 VGND.n90 0.13022
R253 VGND.n92 VGND.n91 0.13022
R254 VGND.n93 VGND.n92 0.13022
R255 VGND.n94 VGND.n93 0.13022
R256 VGND.n95 VGND.n94 0.13022
R257 VGND.n96 VGND.n95 0.13022
R258 VGND.n97 VGND.n96 0.13022
R259 VGND.n98 VGND.n97 0.13022
R260 VGND.n99 VGND.n98 0.13022
R261 VGND.n100 VGND.n99 0.13022
R262 VGND.n101 VGND.n100 0.1133
R263 VGND.n101 VGND.n5 0.07664
R264 VGND.n103 VGND.t5 0.0297714
R265 VGND.n103 VGND.n102 0.0164673
R266 VGND.n106 VGND.n103 0.0164673
R267 VGND.n105 VGND 0.0130333
R268 ua[0].n11 ua[0].n10 8605.04
R269 ua[0].n8 ua[0].n5 8605.04
R270 ua[0].n5 ua[0].n4 3489.23
R271 ua[0].n10 ua[0].n9 3489.23
R272 ua[0].n12 ua[0].n3 1652.71
R273 ua[0].n7 ua[0].n3 1652.71
R274 ua[0].n13 ua[0].n12 1525.46
R275 ua[0].n7 ua[0].n6 1525.46
R276 ua[0].n0 ua[0].t1 660.448
R277 ua[0].n1 ua[0].t3 660.24
R278 ua[0].n13 ua[0].n2 127.248
R279 ua[0].n6 ua[0].n2 127.248
R280 ua[0].n5 ua[0].n2 37.0005
R281 ua[0].n10 ua[0].n3 37.0005
R282 ua[0].n0 ua[0].t0 13.0329
R283 ua[0].n6 ua[0].n1 9.98434
R284 ua[0].n14 ua[0].n13 9.3005
R285 ua[0] ua[0].n15 6.46994
R286 ua[0].n12 ua[0].n11 1.54217
R287 ua[0].n8 ua[0].n7 1.54217
R288 ua[0].n15 ua[0].n0 1.08544
R289 ua[0].n11 ua[0].n4 0.917376
R290 ua[0].n9 ua[0].n8 0.917376
R291 ua[0].n15 ua[0].n14 0.899115
R292 ua[0].n14 ua[0].n1 0.684342
R293 ua[0].n9 ua[0].t2 0.626126
R294 ua[0].t2 ua[0].n4 0.626126
R295 stage1.n9 stage1.n2 741
R296 stage1.n6 stage1.n2 741
R297 stage1.n7 stage1.n6 741
R298 stage1.n5 stage1.t0 323.575
R299 stage1.n9 stage1.n8 236.839
R300 stage1.n5 stage1.n4 151.427
R301 stage1.n3 stage1.n0 146.447
R302 stage1.n3 stage1.n1 146.447
R303 stage1.n10 stage1.n1 139.639
R304 stage1.n11 stage1.n0 133.804
R305 stage1 stage1.t1 69.0795
R306 stage1.n10 stage1.n9 46.2505
R307 stage1.n6 stage1.n3 46.2505
R308 stage1.n6 stage1.n5 46.2505
R309 stage1.n7 stage1.n1 46.2505
R310 stage1.n2 stage1.n0 46.2505
R311 stage1.t0 stage1.n2 46.2505
R312 stage1.n8 stage1.n7 29.6199
R313 stage1.n8 stage1.t0 14.7834
R314 stage1.n12 stage1.n11 5.56832
R315 stage1.n11 stage1.n10 3.2005
R316 stage1 stage1.n12 3.063
R317 stage1.n12 stage1.t2 1.84196
R318 stage2.n9 stage2.n2 741
R319 stage2.n6 stage2.n2 741
R320 stage2.n7 stage2.n6 741
R321 stage2.n5 stage2.t0 323.575
R322 stage2.n9 stage2.n8 236.839
R323 stage2.n5 stage2.n4 151.427
R324 stage2.n3 stage2.n0 146.447
R325 stage2.n3 stage2.n1 146.447
R326 stage2.n10 stage2.n1 132.846
R327 stage2.n11 stage2.n0 129.567
R328 stage2 stage2.t1 69.7157
R329 stage2.n10 stage2.n9 46.2505
R330 stage2.n6 stage2.n3 46.2505
R331 stage2.n6 stage2.n5 46.2505
R332 stage2.n7 stage2.n1 46.2505
R333 stage2.n2 stage2.n0 46.2505
R334 stage2.t0 stage2.n2 46.2505
R335 stage2.n8 stage2.n7 29.6199
R336 stage2.n8 stage2.t0 14.7834
R337 stage2.n12 stage2.n11 5.52342
R338 stage2 stage2.n12 2.89633
R339 stage2.n12 stage2.t2 1.83674
R340 stage2.n11 stage2.n10 1.23921
R341 clk.n0 clk.t1 265.868
R342 clk.n0 clk.t0 236.738
R343 clk.n1 clk.n0 16.0872
R344 clk clk.n1 0.0952833
R345 clk.n1 clk 0.0189314
R346 clka.n0 clka.t1 19.2376
R347 clka.n0 clka.t0 10.2333
R348 clka clka.n0 5.69842
R349 clkb clkb.t2 167.837
R350 clkb clkb.t1 82.955
R351 clkb clkb.t0 9.29528
R352 VAPWR.n9 VAPWR.n3 1053.52
R353 VAPWR.n9 VAPWR.n4 1053.52
R354 VAPWR.n18 VAPWR.n4 1053.52
R355 VAPWR.n18 VAPWR.n3 1053.52
R356 VAPWR.n11 VAPWR.n5 1053.52
R357 VAPWR.n11 VAPWR.n6 1053.52
R358 VAPWR.n16 VAPWR.n6 1053.52
R359 VAPWR.n16 VAPWR.n5 1053.52
R360 VAPWR.n8 VAPWR.n1 206.306
R361 VAPWR.n8 VAPWR.n2 206.306
R362 VAPWR.n12 VAPWR.n7 206.306
R363 VAPWR.n13 VAPWR.n12 206.306
R364 VAPWR.n19 VAPWR.n2 200.638
R365 VAPWR.n15 VAPWR.n7 200.596
R366 VAPWR.n14 VAPWR.n13 200.2
R367 VAPWR.n20 VAPWR.n1 199.446
R368 VAPWR.n0 VAPWR.t1 167.04
R369 VAPWR.n22 VAPWR.t2 167.038
R370 VAPWR.n17 VAPWR.t0 117.51
R371 VAPWR.n10 VAPWR.t0 117.51
R372 VAPWR.n23 VAPWR.t3 71.4739
R373 VAPWR.n3 VAPWR.n1 46.2505
R374 VAPWR.t0 VAPWR.n3 46.2505
R375 VAPWR.n4 VAPWR.n2 46.2505
R376 VAPWR.t0 VAPWR.n4 46.2505
R377 VAPWR.n7 VAPWR.n5 46.2505
R378 VAPWR.n5 VAPWR.t0 46.2505
R379 VAPWR.n13 VAPWR.n6 46.2505
R380 VAPWR.n6 VAPWR.t0 46.2505
R381 VAPWR.n19 VAPWR.n18 23.1255
R382 VAPWR.n18 VAPWR.n17 23.1255
R383 VAPWR.n9 VAPWR.n8 23.1255
R384 VAPWR.n10 VAPWR.n9 23.1255
R385 VAPWR.n12 VAPWR.n11 23.1255
R386 VAPWR.n11 VAPWR.n10 23.1255
R387 VAPWR.n16 VAPWR.n15 23.1255
R388 VAPWR.n17 VAPWR.n16 23.1255
R389 VAPWR.n23 VAPWR.n22 9.14026
R390 VAPWR VAPWR.n23 7.20367
R391 VAPWR.n14 VAPWR.n0 1.163
R392 VAPWR.n21 VAPWR.n20 1.163
R393 VAPWR.n20 VAPWR.n19 1.06717
R394 VAPWR.n21 VAPWR.n0 0.606832
R395 VAPWR.n15 VAPWR.n14 0.356056
R396 VAPWR.n22 VAPWR.n21 0.00251613
C0 VAPWR rst_n 1.03e-19
C1 uio_in[4] uio_in[3] 0.031023f
C2 ui_in[7] ui_in[6] 0.031023f
C3 stage2 stage3 1.1489f
C4 VDPWR m2_2064_15598# 0.294528f
C5 vout VAPWR 0.553317f
C6 ui_in[2] ui_in[1] 0.031023f
C7 VDPWR m2_1280_33406# 0.024041f
C8 VDPWR m2_1056_29654# 0.0364f
C9 clk VAPWR 0.458284f
C10 VAPWR ui_in[6] 1.03e-19
C11 m2_1056_29654# m2_2064_27358# 0.091013f
C12 clkb VAPWR 1.73709f
C13 clk ena 0.034743f
C14 VAPWR stage1 0.51574f
C15 vout ua[0] 0.16305f
C16 ui_in[5] VAPWR 1.03e-19
C17 clkb stage2 57.2718f
C18 clka VAPWR 4.91567f
C19 stage2 stage1 1.20983f
C20 VDPWR m2_2064_35982# 0.030818f
C21 vout stage3 0.416737f
C22 m2_1336_8934# m2_944_13022# 0.017782f
C23 VDPWR m2_2120_12070# 0.0364f
C24 clk ui_in[1] 2.07e-20
C25 uio_in[2] uio_in[1] 0.031023f
C26 VDPWR m2_2064_4230# 0.018568f
C27 clka stage2 0.216306f
C28 VDPWR m2_1336_23326# 0.01539f
C29 VDPWR m2_1056_17838# 0.0208f
C30 m2_2064_35982# m2_2064_39062# 0.162853f
C31 clk rst_n 0.031944f
C32 uio_in[6] uio_in[7] 0.031023f
C33 clkb stage3 0.080496f
C34 m2_1336_23326# m2_2064_27358# 0.138713f
C35 uio_in[6] uio_in[5] 0.031023f
C36 m2_1336_8934# m2_2120_12070# 0.135204f
C37 ui_in[3] VAPWR 1.03e-19
C38 ui_in[5] ui_in[4] 0.031023f
C39 m2_2064_4230# m2_272_4342# 0.559432f
C40 clka stage3 57.1062f
C41 uio_in[2] VAPWR 1.03e-19
C42 clka rst_n 3.03e-19
C43 VAPWR uio_in[1] 1.03e-19
C44 ui_in[0] VAPWR 1.03e-19
C45 uio_in[4] uio_in[5] 0.031023f
C46 ui_in[7] VAPWR 1.03e-19
C47 VDPWR m2_2064_27358# 0.02539f
C48 clka vout 0.021853f
C49 VDPWR m2_2064_42086# 0.029183f
C50 ui_in[2] ui_in[3] 0.031023f
C51 VDPWR m2_2064_39062# 0.297004f
C52 m2_1056_29654# m2_1280_33406# 0.041637f
C53 uio_in[2] uio_in[3] 0.031023f
C54 ui_in[5] ui_in[6] 0.031023f
C55 VDPWR m2_1336_8934# 0.0208f
C56 clka clk 0.371694f
C57 VDPWR m2_272_4342# 1.11311f
C58 clkb stage1 0.165327f
C59 ui_in[3] ui_in[4] 0.031023f
C60 m2_2064_42086# m2_2064_39062# 0.130452f
C61 ui_in[0] ui_in[1] 0.031023f
C62 clka clkb 2.8393f
C63 uio_in[0] uio_in[1] 0.031023f
C64 clka stage1 57.232803f
C65 m2_2064_15598# m2_2120_12070# 0.104769f
C66 ua[1] ua[0] 0.001614f
C67 ui_in[7] uio_in[0] 0.031023f
C68 ui_in[0] rst_n 0.031023f
C69 m2_1336_8934# m2_272_4342# 0.00172f
C70 m2_2064_35982# m2_1280_33406# 0.0711f
C71 m2_2064_15598# m2_1056_17838# 0.151985f
C72 VAPWR uio_in[3] 1.03e-19
C73 VAPWR ua[0] 0.262061f
C74 ui_in[2] VAPWR 1.03e-19
C75 VAPWR ui_in[1] 1.03e-19
C76 VAPWR uio_in[0] 1.03e-19
C77 m2_2120_12070# m2_944_13022# 0.105624f
C78 ui_in[4] VAPWR 1.03e-19
C79 ui_in[0] clk 9.82e-20
C80 ua[1] VGND 0.145965f
C81 ua[2] VGND 0.148302f
C82 ua[3] VGND 0.148302f
C83 ua[4] VGND 0.148302f
C84 ua[5] VGND 0.148302f
C85 ua[6] VGND 0.146962f
C86 ua[7] VGND 0.146962f
C87 VDPWR VGND 20.8487f
C88 ena VGND 0.075936f
C89 rst_n VGND 0.04853f
C90 ui_in[0] VGND 0.048746f
C91 ui_in[1] VGND 0.048746f
C92 ui_in[2] VGND 0.048746f
C93 ui_in[3] VGND 0.048746f
C94 ui_in[4] VGND 0.048746f
C95 ui_in[5] VGND 0.048746f
C96 ui_in[6] VGND 0.048746f
C97 ui_in[7] VGND 0.048746f
C98 uio_in[0] VGND 0.048746f
C99 uio_in[1] VGND 0.048746f
C100 uio_in[2] VGND 0.048746f
C101 uio_in[3] VGND 0.048746f
C102 uio_in[4] VGND 0.048746f
C103 uio_in[5] VGND 0.048746f
C104 uio_in[6] VGND 0.048746f
C105 uio_in[7] VGND 0.079769f
C106 clk VGND 1.74178f
C107 ua[0] VGND 44.30256f
C108 VAPWR VGND 26.80059f
C109 m2_2064_4230# VGND 2.41736f $ **FLOATING
C110 m2_272_4342# VGND 11.7441f $ **FLOATING
C111 m2_1336_8934# VGND 5.1283f $ **FLOATING
C112 m2_2120_12070# VGND 3.18023f $ **FLOATING
C113 m2_944_13022# VGND 0.831538f $ **FLOATING
C114 m2_2064_15598# VGND 5.96367f $ **FLOATING
C115 m2_1056_17838# VGND 4.71527f $ **FLOATING
C116 m2_1336_23326# VGND 4.89346f $ **FLOATING
C117 m2_2064_27358# VGND 4.41841f $ **FLOATING
C118 m2_1056_29654# VGND 4.17312f $ **FLOATING
C119 m2_1280_33406# VGND 4.18017f $ **FLOATING
C120 m2_2064_35982# VGND 4.2612f $ **FLOATING
C121 m2_2064_39062# VGND 5.97958f $ **FLOATING
C122 m2_2064_42086# VGND 4.35936f $ **FLOATING
C123 clkb VGND 17.05209f
C124 clka VGND 32.70971f
C125 vout VGND 0.126327p
C126 stage3 VGND 6.408846f
C127 stage2 VGND 6.986602f
C128 stage1 VGND 7.681975f
C129 VAPWR.t1 VGND 0.004715f
C130 VAPWR.n0 VGND 0.024338f
C131 VAPWR.n1 VGND 0.005645f
C132 VAPWR.n2 VGND 0.005659f
C133 VAPWR.n3 VGND 0.009696f
C134 VAPWR.n4 VGND 0.009696f
C135 VAPWR.t0 VGND 0.107388f
C136 VAPWR.n5 VGND 0.009696f
C137 VAPWR.n6 VGND 0.009696f
C138 VAPWR.n7 VGND 0.00566f
C139 VAPWR.n8 VGND 0.005587f
C140 VAPWR.n9 VGND 0.009493f
C141 VAPWR.n10 VGND 0.10159f
C142 VAPWR.n11 VGND 0.009493f
C143 VAPWR.n12 VGND 0.005587f
C144 VAPWR.n13 VGND 0.005655f
C145 VAPWR.n14 VGND 0.002956f
C146 VAPWR.n15 VGND 0.002961f
C147 VAPWR.n16 VGND 0.009493f
C148 VAPWR.n17 VGND 0.10159f
C149 VAPWR.n18 VGND 0.009493f
C150 VAPWR.n19 VGND 0.002971f
C151 VAPWR.n20 VGND 0.002956f
C152 VAPWR.n21 VGND 0.020654f
C153 VAPWR.t2 VGND 0.004715f
C154 VAPWR.n22 VGND 0.024607f
C155 VAPWR.t3 VGND 0.020636f
C156 VAPWR.n23 VGND 2.35518f
C157 clkb.t0 VGND 58.5911f
C158 clkb.t1 VGND 0.021049f
C159 clkb.t2 VGND 0.033105f
C160 clka.t1 VGND 59.9238f
C161 clka.t0 VGND 58.5954f
C162 clka.n0 VGND 2.92777f
C163 stage2.t2 VGND 55.0583f
C164 stage2.n0 VGND 0.014797f
C165 stage2.n1 VGND 0.014928f
C166 stage2.n2 VGND 0.026188f
C167 stage2.t0 VGND 0.151672f
C168 stage2.n3 VGND 0.015465f
C169 stage2.n4 VGND 0.031658f
C170 stage2.n5 VGND 0.099305f
C171 stage2.n6 VGND 0.026477f
C172 stage2.n7 VGND 0.026188f
C173 stage2.n9 VGND 0.141061f
C174 stage2.n10 VGND 0.010925f
C175 stage2.n11 VGND 0.02724f
C176 stage2.n12 VGND 0.690044f
C177 stage2.t1 VGND 0.052779f
C178 stage1.t2 VGND 54.924603f
C179 stage1.n0 VGND 0.014847f
C180 stage1.n1 VGND 0.015108f
C181 stage1.n2 VGND 0.026122f
C182 stage1.t0 VGND 0.151293f
C183 stage1.n3 VGND 0.015426f
C184 stage1.n4 VGND 0.031578f
C185 stage1.n5 VGND 0.099057f
C186 stage1.n6 VGND 0.026411f
C187 stage1.n7 VGND 0.026122f
C188 stage1.n9 VGND 0.140709f
C189 stage1.n10 VGND 0.009264f
C190 stage1.n11 VGND 0.024349f
C191 stage1.n12 VGND 0.705173f
C192 stage1.t1 VGND 0.052067f
C193 ua[0].t1 VGND 0.005519f
C194 ua[0].t0 VGND 3.10314f
C195 ua[0].n0 VGND 0.276422f
C196 ua[0].t3 VGND 0.005516f
C197 ua[0].n1 VGND 0.026563f
C198 ua[0].n2 VGND 0.014389f
C199 ua[0].n3 VGND 0.182239f
C200 ua[0].n5 VGND 2.08895f
C201 ua[0].n6 VGND 0.091492f
C202 ua[0].n7 VGND 0.173982f
C203 ua[0].n8 VGND 0.307968f
C204 ua[0].t2 VGND 3.44356f
C205 ua[0].n10 VGND 2.08895f
C206 ua[0].n11 VGND 0.307968f
C207 ua[0].n12 VGND 0.173982f
C208 ua[0].n13 VGND 0.090925f
C209 ua[0].n14 VGND 0.014867f
C210 ua[0].n15 VGND 0.090214f
C211 stage3.t1 VGND 0.051318f
C212 stage3.t2 VGND 55.3166f
C213 stage3.n0 VGND 0.015024f
C214 stage3.n1 VGND 0.01533f
C215 stage3.n2 VGND 0.026303f
C216 stage3.t0 VGND 0.152337f
C217 stage3.n3 VGND 0.015532f
C218 stage3.n4 VGND 0.031796f
C219 stage3.n5 VGND 0.09974f
C220 stage3.n6 VGND 0.026593f
C221 stage3.n7 VGND 0.026303f
C222 stage3.n9 VGND 0.14168f
C223 stage3.n10 VGND 0.008747f
C224 stage3.n11 VGND 0.046769f
C225 stage3.n12 VGND 0.429482f
C226 stage3.n13 VGND 0.266759f
C227 vout.t1 VGND 8.153561f
C228 vout.n0 VGND 0.003407f
C229 vout.n1 VGND 0.003437f
C230 vout.n2 VGND 0.005855f
C231 vout.n3 VGND 0.005855f
C232 vout.n4 VGND 0.003458f
C233 vout.n5 VGND 0.031538f
C234 vout.t0 VGND 0.033911f
C235 vout.n7 VGND 0.007078f
C236 vout.n8 VGND 0.022202f
C237 vout.n9 VGND 0.00592f
C238 vout.n10 VGND 0.002234f
C239 vout.n11 VGND 0.080577f
C240 vout.n12 VGND 0.915113f
C241 vout.t3 VGND 0.001141f
C242 vout.n13 VGND 0.020912f
C243 vout.n14 VGND 0.037591f
C244 vout.n15 VGND 0.430897f
C245 vout.n16 VGND 0.430897f
C246 vout.n17 VGND 0.037332f
C247 vout.n18 VGND 0.063526f
C248 vout.t2 VGND 0.71032f
C249 vout.n21 VGND 0.063526f
C250 vout.n22 VGND 0.035065f
C251 vout.n23 VGND 0.02036f
C252 vout.n24 VGND 0.654245f
C253 w_20072_2496.t0 VGND 13.4908f
C254 w_20072_2496.t2 VGND 12.7878f
C255 w_20072_2496.t3 VGND 0.010686f
C256 w_20072_2496.t1 VGND 0.010683f
.ends

