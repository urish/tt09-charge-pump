magic
tech sky130A
magscale 1 2
timestamp 1725639464
<< locali >>
rect 31012 43728 31070 43762
<< viali >>
rect 30512 44468 30570 44502
rect 31012 44466 31070 44500
rect 30336 44280 30370 44340
rect 31212 44302 31246 44356
rect 30336 43620 30370 43680
rect 31212 43542 31246 43596
rect 21184 41780 21322 42604
rect 21836 42124 21884 42272
rect 21184 36156 21322 36980
rect 21842 36484 21904 36656
rect 21188 30744 21326 31568
rect 21844 31082 21884 31260
rect 21316 28248 22008 28342
rect 21424 27664 21484 28092
rect 23276 2902 23312 2948
rect 31490 1966 31530 2000
rect 31490 1478 31530 1512
<< metal1 >>
rect 30500 44502 30760 44520
rect 30500 44468 30512 44502
rect 30570 44468 30760 44502
rect 30500 44460 30760 44468
rect 30820 44506 31080 44520
rect 30820 44500 31082 44506
rect 30820 44466 31012 44500
rect 31070 44466 31082 44500
rect 30820 44460 31082 44466
rect 31200 44360 31260 44520
rect 30330 44340 30376 44352
rect 29150 44280 29160 44340
rect 29340 44280 30336 44340
rect 30370 44280 30480 44340
rect 30580 44300 31000 44360
rect 31100 44356 31260 44360
rect 31100 44302 31212 44356
rect 31246 44302 31260 44356
rect 31100 44300 31260 44302
rect 30330 44268 30376 44280
rect 30760 43980 30820 44300
rect 30750 43920 30760 43980
rect 30820 43920 30830 43980
rect 30760 43780 30820 43920
rect 30480 43720 31100 43780
rect 30330 43680 30376 43692
rect 29150 43620 29160 43680
rect 29340 43620 30336 43680
rect 30370 43620 30480 43680
rect 30330 43608 30376 43620
rect 31200 43600 31260 44300
rect 30600 43540 30980 43600
rect 31100 43596 31260 43600
rect 31100 43542 31212 43596
rect 31246 43542 31260 43596
rect 31100 43540 31260 43542
rect 30680 43140 30740 43540
rect 31200 43400 31260 43540
rect 31190 43280 31200 43400
rect 31260 43280 31270 43400
rect 30650 42960 30660 43140
rect 30780 42960 30790 43140
rect 21178 42604 21328 42616
rect 21174 41780 21184 42604
rect 21322 41780 21332 42604
rect 21830 42274 21890 42284
rect 22166 42274 22320 42300
rect 21560 42104 21570 42274
rect 21740 42104 21750 42274
rect 21830 42272 22320 42274
rect 21830 42124 21836 42272
rect 21884 42124 22320 42272
rect 21830 42120 22320 42124
rect 22500 42120 22510 42300
rect 21830 42112 21890 42120
rect 21178 41768 21328 41780
rect 21178 36980 21328 36992
rect 21174 36156 21184 36980
rect 21322 36156 21332 36980
rect 21836 36660 21910 36668
rect 21836 36656 22320 36660
rect 21568 36476 21578 36656
rect 21758 36476 21768 36656
rect 21836 36484 21842 36656
rect 21904 36484 22320 36656
rect 21836 36480 22320 36484
rect 22500 36480 22510 36660
rect 21836 36472 21910 36480
rect 21178 36144 21328 36156
rect 21182 31568 21332 31580
rect 21178 30744 21188 31568
rect 21326 30744 21336 31568
rect 21838 31260 21890 31272
rect 21560 31074 21570 31246
rect 21742 31074 21752 31246
rect 21838 31082 21844 31260
rect 21884 31242 22514 31260
rect 21884 31096 22362 31242
rect 22498 31096 22514 31242
rect 21884 31082 22514 31096
rect 21838 31080 22514 31082
rect 21838 31070 21890 31080
rect 21182 30732 21332 30744
rect 21144 28354 22128 28356
rect 21142 28226 21152 28354
rect 21336 28342 22128 28354
rect 22008 28248 22128 28342
rect 21336 28226 22128 28248
rect 21144 28212 22128 28226
rect 19380 28146 20220 28200
rect 19380 28140 21496 28146
rect 19370 27900 19380 28140
rect 19620 28092 21496 28140
rect 19620 27900 21424 28092
rect 19380 27664 21424 27900
rect 21484 27664 21496 28092
rect 21558 27786 21568 27966
rect 21748 27786 21758 27966
rect 19380 27660 21496 27664
rect 19370 27420 19380 27660
rect 19620 27610 21496 27660
rect 19620 27420 20220 27610
rect 19380 27180 20220 27420
rect 19370 26940 19380 27180
rect 19620 26940 20220 27180
rect 19380 26880 20220 26940
rect 23060 2898 23070 2960
rect 23126 2948 23136 2960
rect 23270 2948 23318 2960
rect 23126 2902 23276 2948
rect 23312 2902 23429 2948
rect 23126 2898 23136 2902
rect 23270 2890 23318 2902
rect 23383 2793 23429 2902
rect 31490 2752 31530 2902
rect 31442 2706 31530 2752
rect 31490 2392 31530 2706
rect 31460 2246 31470 2392
rect 31538 2246 31548 2392
rect 31490 2006 31530 2246
rect 31478 2000 31542 2006
rect 31478 1966 31490 2000
rect 31530 1966 31542 2000
rect 31478 1960 31542 1966
rect 23394 1132 23496 1864
rect 31490 1518 31530 1960
rect 31478 1512 31542 1518
rect 31478 1478 31490 1512
rect 31530 1478 31542 1512
rect 31478 1472 31542 1478
rect 23394 1032 23404 1132
rect 23488 1032 23498 1132
rect 23394 1020 23496 1032
<< via1 >>
rect 30760 44460 30820 44520
rect 29160 44280 29340 44340
rect 30760 43920 30820 43980
rect 29160 43620 29340 43680
rect 31200 43280 31260 43400
rect 30660 42960 30780 43140
rect 21184 41780 21322 42604
rect 21570 42104 21740 42274
rect 22320 42120 22500 42300
rect 21184 36156 21322 36980
rect 21578 36476 21758 36656
rect 22320 36480 22500 36660
rect 21188 30744 21326 31568
rect 21570 31074 21742 31246
rect 22362 31096 22498 31242
rect 21152 28342 21336 28354
rect 21152 28248 21316 28342
rect 21316 28248 21336 28342
rect 21152 28226 21336 28248
rect 19380 27900 19620 28140
rect 21568 27786 21748 27966
rect 19380 27420 19620 27660
rect 19380 26940 19620 27180
rect 23070 2898 23126 2960
rect 31470 2246 31538 2392
rect 23404 1032 23488 1132
<< metal2 >>
rect 28750 45042 28850 45052
rect 28750 44932 28850 44942
rect 28770 44882 28830 44932
rect 28770 44822 30820 44882
rect 30760 44520 30820 44822
rect 30760 44450 30820 44460
rect 29160 44340 29340 44350
rect 29160 44270 29340 44280
rect 27900 43980 28020 43990
rect 30760 43980 30820 43990
rect 28020 43920 30760 43980
rect 30820 43920 30840 43980
rect 28020 43860 30840 43920
rect 27900 43850 28020 43860
rect 29160 43680 29340 43690
rect 29160 43610 29340 43620
rect 21184 42604 21322 42614
rect 22320 42300 22500 42310
rect 21570 42274 21740 42284
rect 21570 42094 21740 42104
rect 21184 41770 21322 41780
rect 22320 37344 22500 42120
rect 21562 37164 22500 37344
rect 21184 36980 21322 36990
rect 21562 36666 21742 37164
rect 21562 36656 21758 36666
rect 21562 36476 21578 36656
rect 21562 36474 21758 36476
rect 21578 36466 21758 36474
rect 22320 36660 22500 36670
rect 21184 36146 21322 36156
rect 22320 32132 22500 36480
rect 21562 31952 22500 32132
rect 29580 32040 29700 43860
rect 31200 43400 31260 43410
rect 31200 43270 31260 43280
rect 30660 43140 30780 43150
rect 30660 42950 30780 42960
rect 21188 31568 21326 31578
rect 21562 31246 21742 31952
rect 29580 31910 29700 31920
rect 21562 31074 21570 31246
rect 21562 31072 21742 31074
rect 21570 31064 21742 31072
rect 22336 31242 22516 31256
rect 22336 31096 22362 31242
rect 22498 31096 22516 31242
rect 21188 30734 21326 30744
rect 22336 28980 22516 31096
rect 21568 28800 22516 28980
rect 21152 28354 21336 28364
rect 21152 28216 21336 28226
rect 19380 28140 19620 28150
rect 19380 27890 19620 27900
rect 21568 27966 21748 28800
rect 21568 27776 21748 27786
rect 19380 27660 19620 27670
rect 19380 27410 19620 27420
rect 19380 27180 19620 27190
rect 19380 26930 19620 26940
rect 23070 2960 23126 2970
rect 23070 2888 23126 2898
rect 31470 2392 31538 2402
rect 31470 2236 31538 2246
rect 9900 1140 10020 1150
rect 23404 1140 23488 1142
rect 10020 1132 23494 1140
rect 10020 1032 23404 1132
rect 23488 1032 23494 1132
rect 10020 1020 23494 1032
rect 9900 1010 10020 1020
<< via2 >>
rect 28750 44942 28850 45042
rect 29160 44280 29340 44340
rect 27900 43860 28020 43980
rect 29160 43620 29340 43680
rect 21184 41780 21322 42604
rect 21570 42104 21740 42274
rect 22320 42120 22500 42300
rect 21184 36156 21322 36980
rect 22320 36480 22500 36660
rect 31200 43280 31260 43400
rect 30660 42960 30780 43140
rect 21188 30744 21326 31568
rect 29580 31920 29700 32040
rect 22362 31096 22498 31242
rect 21152 28226 21336 28354
rect 19380 27900 19620 28140
rect 19380 27420 19620 27660
rect 19380 26940 19620 27180
rect 23070 2898 23126 2960
rect 31470 2246 31538 2392
rect 9900 1020 10020 1140
<< metal3 >>
rect 28740 45042 28860 45047
rect 28740 44942 28750 45042
rect 28850 44942 28860 45042
rect 28740 44937 28860 44942
rect 29090 44500 29100 44700
rect 29400 44500 29410 44700
rect 29100 44340 29400 44500
rect 29100 44280 29160 44340
rect 29340 44280 29400 44340
rect 27890 43980 28030 43985
rect 27890 43860 27900 43980
rect 28020 43860 28030 43980
rect 27890 43855 28030 43860
rect 29100 43680 29400 44280
rect 21560 43500 28640 43680
rect 29100 43620 29160 43680
rect 29340 43620 29400 43680
rect 29100 43600 29400 43620
rect 21174 42604 21332 42609
rect 21174 41780 21184 42604
rect 21322 41780 21332 42604
rect 21560 42279 21740 43500
rect 28460 43440 28640 43500
rect 28432 43260 28440 43440
rect 28740 43400 28750 43440
rect 31190 43400 31270 43405
rect 28740 43280 31200 43400
rect 31260 43280 31270 43400
rect 28740 43260 28750 43280
rect 31190 43275 31270 43280
rect 28460 43246 28640 43260
rect 30650 43140 30790 43145
rect 30650 42960 30660 43140
rect 30780 42960 30790 43140
rect 30650 42955 30790 42960
rect 22310 42300 22510 42305
rect 21560 42274 21750 42279
rect 21560 42104 21570 42274
rect 21740 42104 21750 42274
rect 22310 42120 22320 42300
rect 22500 42120 22510 42300
rect 22310 42115 22510 42120
rect 21560 42099 21750 42104
rect 21560 42088 21740 42099
rect 21174 41775 21332 41780
rect 30660 37440 30780 42955
rect 28070 37320 28080 37440
rect 28260 37320 30780 37440
rect 21174 36980 21332 36985
rect 21174 36156 21184 36980
rect 21322 36156 21332 36980
rect 22310 36660 22510 36665
rect 22310 36480 22320 36660
rect 22500 36480 22510 36660
rect 22310 36475 22510 36480
rect 21174 36151 21332 36156
rect 29570 32040 29710 32045
rect 28070 31920 28080 32040
rect 28260 31920 29580 32040
rect 29700 31920 29710 32040
rect 29570 31915 29710 31920
rect 21178 31568 21336 31573
rect 21178 30744 21188 31568
rect 21326 30744 21336 31568
rect 22352 31242 22508 31247
rect 22352 31096 22362 31242
rect 22498 31096 22508 31242
rect 22352 31091 22508 31096
rect 21178 30739 21336 30744
rect 21142 28354 21346 28359
rect 21142 28226 21152 28354
rect 21336 28226 21346 28354
rect 21142 28221 21346 28226
rect 19380 28145 19620 28200
rect 19370 28140 19630 28145
rect 19370 27900 19380 28140
rect 19620 27900 19630 28140
rect 19370 27895 19630 27900
rect 19380 27665 19620 27895
rect 19370 27660 19630 27665
rect 19370 27420 19380 27660
rect 19620 27420 19630 27660
rect 19370 27415 19630 27420
rect 19380 27185 19620 27415
rect 19370 27180 19630 27185
rect 19370 26940 19380 27180
rect 19620 26940 19630 27180
rect 19370 26935 19630 26940
rect 19380 3136 19620 26935
rect 19380 2965 23130 3136
rect 19380 2960 23136 2965
rect 19380 2898 23070 2960
rect 23126 2898 23136 2960
rect 19380 2896 23136 2898
rect 23060 2893 23136 2896
rect 31460 2392 31548 2397
rect 31460 2246 31470 2392
rect 31538 2246 31548 2392
rect 31460 2241 31548 2246
rect 9890 1140 10030 1145
rect 9890 1020 9900 1140
rect 10020 1020 10030 1140
rect 9890 1015 10030 1020
<< via3 >>
rect 28750 44942 28850 45042
rect 29100 44500 29400 44700
rect 27900 43860 28020 43980
rect 21184 41780 21322 42604
rect 28440 43260 28740 43440
rect 22320 42120 22500 42300
rect 28080 37320 28260 37440
rect 21184 36156 21322 36980
rect 22320 36480 22500 36660
rect 28080 31920 28260 32040
rect 21188 30744 21326 31568
rect 22362 31096 22498 31242
rect 21152 28226 21336 28354
rect 19380 27900 19620 28140
rect 19380 27420 19620 27660
rect 19380 26940 19620 27180
rect 31470 2246 31538 2392
rect 9900 1020 10020 1140
<< metal4 >>
rect 6134 44700 6194 45152
rect 6686 44700 6746 45152
rect 7238 44700 7298 45152
rect 7790 44700 7850 45152
rect 8342 44700 8402 45152
rect 8894 44700 8954 45152
rect 9446 44700 9506 45152
rect 9998 44700 10058 45152
rect 10550 44700 10610 45152
rect 11102 44700 11162 45152
rect 11654 44700 11714 45152
rect 12206 44700 12266 45152
rect 12758 44700 12818 45152
rect 13310 44700 13370 45152
rect 13862 44700 13922 45152
rect 14414 44700 14474 45152
rect 14966 44700 15026 45152
rect 15518 44700 15578 45152
rect 16070 44700 16130 45152
rect 16622 44700 16682 45152
rect 17174 44700 17234 45152
rect 17726 44700 17786 45152
rect 18278 44700 18338 45152
rect 18830 44700 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 45043 28826 45152
rect 28749 45042 28851 45043
rect 28749 44942 28750 45042
rect 28850 44942 28851 45042
rect 29318 44952 29378 45152
rect 28749 44941 28851 44942
rect 29099 44700 29401 44701
rect 6126 44500 29100 44700
rect 29400 44500 29401 44700
rect 9800 27840 10100 44500
rect 21146 42604 21346 44500
rect 29099 44499 29401 44500
rect 27899 43980 28021 43981
rect 27899 43860 27900 43980
rect 28020 43860 28021 43980
rect 27899 43859 28021 43860
rect 27900 43020 28020 43859
rect 28440 43441 28740 44152
rect 28439 43440 28741 43441
rect 28439 43260 28440 43440
rect 28740 43260 28741 43440
rect 28439 43259 28741 43260
rect 21146 41780 21184 42604
rect 21322 41780 21346 42604
rect 22319 42300 22501 42301
rect 22319 42120 22320 42300
rect 22500 42120 22920 42300
rect 22319 42119 22501 42120
rect 21146 36980 21346 41780
rect 27900 37440 28320 37620
rect 27900 37320 28080 37440
rect 28260 37320 28320 37440
rect 27900 37200 28320 37320
rect 21146 36156 21184 36980
rect 21322 36156 21346 36980
rect 22319 36660 22501 36661
rect 22319 36480 22320 36660
rect 22500 36480 22860 36660
rect 22319 36479 22501 36480
rect 21146 31568 21346 36156
rect 27900 32040 28320 32160
rect 27900 31920 28080 32040
rect 28260 31920 28320 32040
rect 27900 31800 28320 31920
rect 21146 30744 21188 31568
rect 21326 30744 21346 31568
rect 22352 31242 22860 31260
rect 22352 31096 22362 31242
rect 22498 31096 22860 31242
rect 22352 31080 22860 31096
rect 21146 28354 21346 30744
rect 21146 28226 21152 28354
rect 21336 28226 21346 28354
rect 21146 28216 21346 28226
rect 19020 28141 19620 28200
rect 19020 28140 19621 28141
rect 19020 27900 19380 28140
rect 19620 27900 19621 28140
rect 19020 27899 19621 27900
rect 9800 25680 13080 27840
rect 19020 27661 19620 27899
rect 19020 27660 19621 27661
rect 19020 27420 19380 27660
rect 19620 27420 19621 27660
rect 19020 27419 19621 27420
rect 19020 27181 19620 27419
rect 19020 27180 19621 27181
rect 19020 26940 19380 27180
rect 19620 26940 19621 27180
rect 19020 26939 19621 26940
rect 19020 26880 19620 26939
rect 9800 1140 10100 25680
rect 9800 1020 9900 1140
rect 10020 1020 10100 1140
rect 9800 1000 10100 1020
rect 28440 1000 28740 43259
rect 31282 2392 31554 2408
rect 31282 2246 31470 2392
rect 31538 2246 31554 2392
rect 31282 2228 31554 2246
rect 31282 780 31462 2228
rect 30362 600 31462 780
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C1
timestamp 1711870259
transform 1 0 25350 0 1 40500
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C2
timestamp 1711870259
transform 1 0 25330 0 1 35060
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C3
timestamp 1711870259
transform 1 0 25330 0 1 29600
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_WMZ6NR  C4
timestamp 1711870259
transform 1 0 15990 0 1 26540
box -3150 -2600 3149 2600
use high_voltage_logo  high_voltage_logo_0
timestamp 1711967973
transform 0 -1 7568 1 0 1262
box 0 0 42336 5768
use sky130_fd_pr__pfet_01v8_BFP3TE  M1
timestamp 1711870259
transform 1 0 31041 0 1 44269
box -241 -369 241 369
use sky130_fd_pr__pfet_01v8_BFP3TE  M2
timestamp 1711870259
transform 1 0 31041 0 1 43531
box -241 -369 241 369
use sky130_fd_pr__nfet_01v8_DSY3K9  M3
timestamp 1711870259
transform -1 0 30541 0 1 44330
box -241 -310 241 310
use sky130_fd_pr__nfet_01v8_DSY3K9  M4
timestamp 1711870259
transform 1 0 30541 0 1 43592
box -241 -310 241 310
use sky130_fd_pr__pfet_g5v0d10v5_RSSSV2  M9
timestamp 1717238374
transform 1 0 27458 0 1 2835
box -4258 -339 4258 339
use sky130_fd_pr__pfet_g5v0d10v5_RSSSV2  M10
timestamp 1717238374
transform 1 0 27458 0 1 1739
box -4258 -339 4258 339
use sky130_fd_pr__diode_pd2nw_11v0_AZAYX8  sky130_fd_pr__diode_pd2nw_11v0_AZAYX8_1
timestamp 1725619700
transform 1 0 21658 0 1 42186
box -478 -478 478 478
use sky130_fd_pr__diode_pd2nw_11v0_AZAYX8  sky130_fd_pr__diode_pd2nw_11v0_AZAYX8_2
timestamp 1725619700
transform 1 0 21666 0 1 36564
box -478 -478 478 478
use sky130_fd_pr__diode_pd2nw_11v0_AZAYX8  sky130_fd_pr__diode_pd2nw_11v0_AZAYX8_3
timestamp 1725619700
transform 1 0 21660 0 1 31156
box -478 -478 478 478
use sky130_fd_pr__diode_pd2nw_11v0_AZAYX8  sky130_fd_pr__diode_pd2nw_11v0_AZAYX8_4
timestamp 1725619700
transform 1 0 21660 0 1 27872
box -478 -478 478 478
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal1 30760 43980 30820 44100 0 FreeSans 320 90 0 0 clka
flabel metal1 30680 42960 30740 43560 0 FreeSans 320 90 0 0 clkb
flabel metal2 22320 37800 22500 42120 0 FreeSans 1600 0 0 0 stage1
flabel metal2 22320 32400 22500 36480 0 FreeSans 1600 0 0 0 stage2
flabel metal3 19380 21660 19620 23880 0 FreeSans 1600 0 0 0 vout
flabel metal2 22336 28800 22516 31080 0 FreeSans 1600 0 0 0 stage3
flabel metal4 28440 1000 28740 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
