* NGSPICE file created from tt_um_urish_charge_pump.ext - technology: sky130A

.subckt tt_um_urish_charge_pump clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VPWR VGND
X0 clka clk.t0 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.45
X1 stage2.t1 clkb.t0 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X2 ua[0].t3 VGND.t3 VGND.t4 ua[0].t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=40
X3 VGND.t5 vout.t2 sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X4 stage3.t1 clka.t1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
D0 stage3.t2 vout.t3 sky130_fd_pr__diode_pd2nw_11v0 pj=4e+06 area=1e+12
X5 clkb.t2 clka VGND.t2 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.45
X6 VPWR.t1 clk.t1 clka VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.45
X7 ua[0].t1 ua[0].t0 vout.t1 vout.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=40
D1 stage1.t1 stage2.t0 sky130_fd_pr__diode_pd2nw_11v0 pj=4e+06 area=1e+12
D2 stage2.t2 stage3.t0 sky130_fd_pr__diode_pd2nw_11v0 pj=4e+06 area=1e+12
D3 VPWR.t3 stage1.t0 sky130_fd_pr__diode_pd2nw_11v0 pj=4e+06 area=1e+12
X8 stage1.t2 clka.t0 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X9 VPWR.t2 clka.t2 clkb.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.45
R0 clk.n0 clk.t1 276.433
R1 clk.n0 clk.t0 244.831
R2 clk.n1 clk.n0 16.3372
R3 clk clk.n1 0.0952833
R4 clk.n1 clk 0.0189314
R5 VGND.n61 VGND.n16 2.0933e+06
R6 VGND.n45 VGND.n18 2.0614e+06
R7 VGND.n51 VGND.n18 1.98293e+06
R8 VGND.n51 VGND.n16 350350
R9 VGND.n62 VGND.n61 196218
R10 VGND.n14 VGND.n11 24077.4
R11 VGND.n52 VGND.n51 18002.7
R12 VGND.n51 VGND.n50 18002.7
R13 VGND.n46 VGND.n45 17143.9
R14 VGND.n45 VGND.n44 17143.9
R15 VGND.n60 VGND.n18 14202.2
R16 VGND.n40 VGND.n39 9131.66
R17 VGND.n39 VGND.n29 9131.66
R18 VGND.n61 VGND.n17 9057.83
R19 VGND.n63 VGND.n62 8780.1
R20 VGND.n30 VGND.n26 7946.72
R21 VGND.n62 VGND.n15 2745.53
R22 VGND.n50 VGND.n19 2624.6
R23 VGND.n46 VGND.n19 2624.6
R24 VGND.n50 VGND.n20 2624.6
R25 VGND.n46 VGND.n20 2624.6
R26 VGND.n33 VGND.n29 2624.6
R27 VGND.n33 VGND.n31 2624.6
R28 VGND.n37 VGND.n31 2624.6
R29 VGND.n37 VGND.n29 2624.6
R30 VGND.n44 VGND.n23 2624.6
R31 VGND.n40 VGND.n23 2624.6
R32 VGND.n44 VGND.n24 2624.6
R33 VGND.n40 VGND.n24 2624.6
R34 VGND.n55 VGND.n17 2624.6
R35 VGND.n55 VGND.n52 2624.6
R36 VGND.n59 VGND.n17 2624.6
R37 VGND.n59 VGND.n52 2624.6
R38 VGND.n13 VGND.n9 2479.88
R39 VGND.n13 VGND.n10 2479.88
R40 VGND.n73 VGND.n9 2479.88
R41 VGND.n73 VGND.n10 2479.88
R42 VGND.n72 VGND.n66 2479.88
R43 VGND.n66 VGND.n64 2479.88
R44 VGND.n65 VGND.n64 2479.88
R45 VGND.n72 VGND.n65 2479.88
R46 VGND.n45 VGND.n22 1219.27
R47 VGND.n28 VGND.n27 1216.4
R48 VGND.n45 VGND.n14 1084.89
R49 VGND.n39 VGND.n22 740.399
R50 VGND.n39 VGND.n38 740.399
R51 VGND.n97 VGND.t4 660.787
R52 VGND.t0 VGND.n11 415.678
R53 VGND.t0 VGND.n63 415.678
R54 VGND.n39 VGND.n28 369.329
R55 VGND.n39 VGND.n26 369.329
R56 VGND.n49 VGND.n21 304.565
R57 VGND.n47 VGND.n21 304.565
R58 VGND.n49 VGND.n48 304.565
R59 VGND.n48 VGND.n47 304.565
R60 VGND.n34 VGND.n32 304.565
R61 VGND.n35 VGND.n34 304.565
R62 VGND.n36 VGND.n35 304.565
R63 VGND.n36 VGND.n32 304.565
R64 VGND.n43 VGND.n42 304.565
R65 VGND.n42 VGND.n41 304.565
R66 VGND.n41 VGND.n25 304.565
R67 VGND.n43 VGND.n25 304.565
R68 VGND.n58 VGND.n53 304.565
R69 VGND.n58 VGND.n57 304.565
R70 VGND.n57 VGND.n56 304.565
R71 VGND.n56 VGND.n53 304.565
R72 VGND.n62 VGND.n14 292.228
R73 VGND.n74 VGND.n73 195
R74 VGND.n73 VGND.t0 195
R75 VGND.n13 VGND.n12 195
R76 VGND.t0 VGND.n13 195
R77 VGND.n72 VGND.n71 195
R78 VGND.t0 VGND.n72 195
R79 VGND.n68 VGND.n64 195
R80 VGND.t0 VGND.n64 195
R81 VGND.n38 VGND.n30 183.243
R82 VGND.n12 VGND.n8 161.13
R83 VGND.n12 VGND.n7 161.13
R84 VGND.n74 VGND.n8 161.13
R85 VGND.n71 VGND.n67 161.13
R86 VGND.n68 VGND.n67 161.13
R87 VGND.n69 VGND.n68 161.13
R88 VGND.n61 VGND.n60 155.025
R89 VGND.n75 VGND.n74 153.601
R90 VGND.n71 VGND.n70 139.294
R91 VGND.n10 VGND.n7 117.001
R92 VGND.n63 VGND.n10 117.001
R93 VGND.n9 VGND.n8 117.001
R94 VGND.n11 VGND.n9 117.001
R95 VGND.n67 VGND.n65 117.001
R96 VGND.n65 VGND.n11 117.001
R97 VGND.n69 VGND.n66 117.001
R98 VGND.n66 VGND.n63 117.001
R99 VGND.n6 VGND.t2 84.0308
R100 VGND.n76 VGND.t1 83.9547
R101 VGND.n54 VGND.n16 68.272
R102 VGND.n32 VGND.n29 58.5005
R103 VGND.n41 VGND.n40 58.5005
R104 VGND.n44 VGND.n43 58.5005
R105 VGND.n47 VGND.n46 58.5005
R106 VGND.n50 VGND.n49 58.5005
R107 VGND.n57 VGND.n52 58.5005
R108 VGND.n53 VGND.n17 58.5005
R109 VGND.n59 VGND.n58 58.5005
R110 VGND.n60 VGND.n59 58.5005
R111 VGND.n34 VGND.n33 58.5005
R112 VGND.n33 VGND.n26 58.5005
R113 VGND.n42 VGND.n24 58.5005
R114 VGND.n28 VGND.n24 58.5005
R115 VGND.n48 VGND.n20 58.5005
R116 VGND.n27 VGND.n20 58.5005
R117 VGND.n35 VGND.n31 58.5005
R118 VGND.n31 VGND.n30 58.5005
R119 VGND.n37 VGND.n36 58.5005
R120 VGND.n38 VGND.n37 58.5005
R121 VGND.n25 VGND.n23 58.5005
R122 VGND.n23 VGND.n22 58.5005
R123 VGND.n21 VGND.n19 58.5005
R124 VGND.n19 VGND.n15 58.5005
R125 VGND.n56 VGND.n55 58.5005
R126 VGND.n55 VGND.n54 58.5005
R127 VGND.n98 VGND.n97 26.0302
R128 VGND.n27 VGND.n18 24.0676
R129 VGND.n70 VGND.n69 21.8358
R130 VGND.n76 VGND.n75 9.3005
R131 VGND.n70 VGND.n6 9.3005
R132 VGND.n75 VGND.n7 7.52991
R133 VGND.n97 VGND.t3 7.28674
R134 VGND.n77 VGND.n6 5.60682
R135 VGND.n77 VGND.n76 5.50342
R136 VGND.n54 VGND.n15 5.10491
R137 VGND.n95 VGND 4.20543
R138 VGND.n99 VGND.n98 3.8545
R139 VGND.n78 VGND.n77 3.05557
R140 VGND.n95 VGND.n94 2.62623
R141 VGND VGND.n99 0.365382
R142 VGND.n0 uio_oe[7] 0.32762
R143 VGND.n94 uio_oe[0] 0.213567
R144 VGND.n78 uo_out[0] 0.1979
R145 VGND.n79 uo_out[1] 0.1979
R146 VGND.n80 uo_out[2] 0.1979
R147 VGND.n81 uo_out[3] 0.1979
R148 VGND.n82 uo_out[4] 0.1979
R149 VGND.n83 uo_out[5] 0.1979
R150 VGND.n84 uo_out[6] 0.1979
R151 VGND.n85 uo_out[7] 0.1979
R152 VGND.n86 uio_out[0] 0.1979
R153 VGND.n87 uio_out[1] 0.1979
R154 VGND.n88 uio_out[2] 0.1979
R155 VGND.n89 uio_out[3] 0.1979
R156 VGND.n90 uio_out[4] 0.1979
R157 VGND.n91 uio_out[5] 0.1979
R158 VGND.n92 uio_out[6] 0.1979
R159 VGND.n93 uio_out[7] 0.1979
R160 VGND.n5 uio_oe[1] 0.1979
R161 VGND.n4 uio_oe[2] 0.1979
R162 VGND.n3 uio_oe[3] 0.1979
R163 VGND.n2 uio_oe[4] 0.1979
R164 VGND.n1 uio_oe[5] 0.1979
R165 VGND.n0 uio_oe[6] 0.1979
R166 VGND.n5 VGND.n4 0.13022
R167 VGND.n4 VGND.n3 0.13022
R168 VGND.n3 VGND.n2 0.13022
R169 VGND.n2 VGND.n1 0.13022
R170 VGND.n1 VGND.n0 0.13022
R171 VGND.n79 VGND.n78 0.13022
R172 VGND.n80 VGND.n79 0.13022
R173 VGND.n81 VGND.n80 0.13022
R174 VGND.n82 VGND.n81 0.13022
R175 VGND.n83 VGND.n82 0.13022
R176 VGND.n84 VGND.n83 0.13022
R177 VGND.n85 VGND.n84 0.13022
R178 VGND.n86 VGND.n85 0.13022
R179 VGND.n87 VGND.n86 0.13022
R180 VGND.n88 VGND.n87 0.13022
R181 VGND.n89 VGND.n88 0.13022
R182 VGND.n90 VGND.n89 0.13022
R183 VGND.n91 VGND.n90 0.13022
R184 VGND.n92 VGND.n91 0.13022
R185 VGND.n93 VGND.n92 0.13022
R186 VGND.n94 VGND.n93 0.1133
R187 VGND.n94 VGND.n5 0.07664
R188 VGND.n96 VGND.t5 0.0297714
R189 VGND.n96 VGND.n95 0.0164673
R190 VGND.n99 VGND.n96 0.0164673
R191 VGND.n98 VGND 0.0130333
R192 clka clka.t2 276.433
R193 clka.n0 clka.t1 19.2376
R194 clka.n0 clka.t0 10.2333
R195 clka clka.n0 6.03696
R196 stage2.n9 stage2.n2 741
R197 stage2.n6 stage2.n2 741
R198 stage2.n7 stage2.n6 741
R199 stage2.n5 stage2.t0 323.575
R200 stage2.n9 stage2.n8 236.839
R201 stage2.n5 stage2.n4 151.427
R202 stage2.n3 stage2.n0 146.447
R203 stage2.n3 stage2.n1 146.447
R204 stage2.n10 stage2.n1 132.846
R205 stage2.n11 stage2.n0 129.567
R206 stage2 stage2.t2 69.7157
R207 stage2.n10 stage2.n9 46.2505
R208 stage2.n6 stage2.n3 46.2505
R209 stage2.n6 stage2.n5 46.2505
R210 stage2.n7 stage2.n1 46.2505
R211 stage2.n2 stage2.n0 46.2505
R212 stage2.t0 stage2.n2 46.2505
R213 stage2.n8 stage2.n7 29.6199
R214 stage2.n8 stage2.t0 14.7834
R215 stage2.n12 stage2.n11 5.52342
R216 stage2 stage2.n12 2.89633
R217 stage2.n12 stage2.t1 1.83674
R218 stage2.n11 stage2.n10 1.23921
R219 clkb clkb.t1 167.643
R220 clkb clkb.t2 83.7335
R221 clkb clkb.t0 9.32862
R222 ua[0].n11 ua[0].n10 8605.04
R223 ua[0].n8 ua[0].n5 8605.04
R224 ua[0].n5 ua[0].n4 3489.23
R225 ua[0].n10 ua[0].n9 3489.23
R226 ua[0].n12 ua[0].n3 1652.71
R227 ua[0].n7 ua[0].n3 1652.71
R228 ua[0].n13 ua[0].n12 1525.46
R229 ua[0].n7 ua[0].n6 1525.46
R230 ua[0].n0 ua[0].t1 660.448
R231 ua[0].n1 ua[0].t3 660.24
R232 ua[0].n13 ua[0].n2 127.248
R233 ua[0].n6 ua[0].n2 127.248
R234 ua[0].n5 ua[0].n2 37.0005
R235 ua[0].n10 ua[0].n3 37.0005
R236 ua[0].n0 ua[0].t0 13.0329
R237 ua[0].n6 ua[0].n1 9.98434
R238 ua[0].n14 ua[0].n13 9.3005
R239 ua[0] ua[0].n15 6.46994
R240 ua[0].n12 ua[0].n11 1.54217
R241 ua[0].n8 ua[0].n7 1.54217
R242 ua[0].n15 ua[0].n0 1.08544
R243 ua[0].n11 ua[0].n4 0.917376
R244 ua[0].n9 ua[0].n8 0.917376
R245 ua[0].n15 ua[0].n14 0.899115
R246 ua[0].n14 ua[0].n1 0.684342
R247 ua[0].n9 ua[0].t2 0.626126
R248 ua[0].t2 ua[0].n4 0.626126
R249 vout.n21 vout.n20 8605.04
R250 vout.n18 vout.n16 8605.04
R251 vout.n21 vout.n15 3489.23
R252 vout.n19 vout.n18 3489.23
R253 vout.n17 vout.n13 1652.71
R254 vout.n17 vout.n14 1652.71
R255 vout.n22 vout.n14 1652.71
R256 vout.n23 vout.n13 1618.34
R257 vout.n5 vout.n2 741
R258 vout.n9 vout.n2 741
R259 vout.n9 vout.n3 741
R260 vout.n24 vout.t1 660.668
R261 vout.n8 vout.t3 323.575
R262 vout.n6 vout.n5 236.839
R263 vout.n8 vout.n7 151.427
R264 vout.n4 vout.n0 146.447
R265 vout.n4 vout.n1 146.447
R266 vout.n10 vout.n1 125.314
R267 vout.n11 vout.n0 123.569
R268 vout.n5 vout.n4 46.2505
R269 vout.n10 vout.n9 46.2505
R270 vout.n9 vout.n8 46.2505
R271 vout.n3 vout.n1 46.2505
R272 vout.n2 vout.n0 46.2505
R273 vout.t3 vout.n2 46.2505
R274 vout.n18 vout.n17 37.0005
R275 vout.n22 vout.n21 37.0005
R276 vout.n23 vout.n22 33.4018
R277 vout.n6 vout.n3 29.6199
R278 vout.t3 vout.n6 14.7834
R279 vout vout.n24 12.7263
R280 vout.n24 vout.n23 9.3005
R281 vout.n12 vout.n11 2.16948
R282 vout.n11 vout.n10 1.74595
R283 vout.n16 vout.n13 1.54217
R284 vout.n20 vout.n14 1.54217
R285 vout vout.n12 1.09447
R286 vout.n16 vout.n15 0.917376
R287 vout.n20 vout.n19 0.917376
R288 vout.n19 vout.t0 0.626126
R289 vout.t0 vout.n15 0.626126
R290 vout.n12 vout.t2 0.404364
R291 stage3.n9 stage3.n2 741
R292 stage3.n6 stage3.n2 741
R293 stage3.n7 stage3.n6 741
R294 stage3.n5 stage3.t0 323.575
R295 stage3.n9 stage3.n8 236.839
R296 stage3.n5 stage3.n4 151.427
R297 stage3.n3 stage3.n0 146.447
R298 stage3.n3 stage3.n1 146.447
R299 stage3.n10 stage3.n1 142.268
R300 stage3.n11 stage3.n0 135.774
R301 stage3 stage3.t2 68.9393
R302 stage3.n10 stage3.n9 46.2505
R303 stage3.n6 stage3.n3 46.2505
R304 stage3.n6 stage3.n5 46.2505
R305 stage3.n7 stage3.n1 46.2505
R306 stage3.n2 stage3.n0 46.2505
R307 stage3.t0 stage3.n2 46.2505
R308 stage3.n8 stage3.n7 29.6199
R309 stage3.n8 stage3.t0 14.7834
R310 stage3.n11 stage3.n10 4.8005
R311 stage3.n12 stage3.n11 4.61856
R312 stage3.n12 stage3.t1 2.68428
R313 stage3.n13 stage3.n12 1.52064
R314 stage3 stage3.n13 0.1255
R315 stage3.n13 stage3 0.063
R316 VPWR.n16 VPWR.n5 1718.82
R317 VPWR.n12 VPWR.n5 1718.82
R318 VPWR.n16 VPWR.n6 1718.82
R319 VPWR.n12 VPWR.n6 1718.82
R320 VPWR.n10 VPWR.n3 1718.82
R321 VPWR.n10 VPWR.n4 1718.82
R322 VPWR.n18 VPWR.n4 1718.82
R323 VPWR.n18 VPWR.n3 1718.82
R324 VPWR.n13 VPWR.n8 183.341
R325 VPWR.n15 VPWR.n14 183.341
R326 VPWR.n14 VPWR.n13 183.341
R327 VPWR.n9 VPWR.n1 183.341
R328 VPWR.n9 VPWR.n2 183.341
R329 VPWR.n19 VPWR.n2 183.341
R330 VPWR.n20 VPWR.n1 169.036
R331 VPWR.n0 VPWR.t1 167.94
R332 VPWR.n21 VPWR.t2 167.881
R333 VPWR.n8 VPWR.n7 160.754
R334 VPWR.n17 VPWR.t0 121.004
R335 VPWR.n11 VPWR.t0 121.004
R336 VPWR.n23 VPWR.t3 71.4739
R337 VPWR.n14 VPWR.n6 61.6672
R338 VPWR.n6 VPWR.t0 61.6672
R339 VPWR.n8 VPWR.n5 61.6672
R340 VPWR.n5 VPWR.t0 61.6672
R341 VPWR.n3 VPWR.n1 61.6672
R342 VPWR.t0 VPWR.n3 61.6672
R343 VPWR.n4 VPWR.n2 61.6672
R344 VPWR.t0 VPWR.n4 61.6672
R345 VPWR.n13 VPWR.n12 26.4291
R346 VPWR.n12 VPWR.n11 26.4291
R347 VPWR.n16 VPWR.n15 26.4291
R348 VPWR.n17 VPWR.n16 26.4291
R349 VPWR.n10 VPWR.n9 26.4291
R350 VPWR.n11 VPWR.n10 26.4291
R351 VPWR.n19 VPWR.n18 26.4291
R352 VPWR.n18 VPWR.n17 26.4291
R353 VPWR.n15 VPWR.n7 22.5887
R354 VPWR.n20 VPWR.n19 14.3064
R355 VPWR.n7 VPWR.n0 9.3005
R356 VPWR.n21 VPWR.n20 9.3005
R357 VPWR VPWR.n23 7.20367
R358 VPWR.n23 VPWR.n22 7.05903
R359 VPWR.n22 VPWR.n0 1.46092
R360 VPWR.n22 VPWR.n21 0.00258333
R361 stage1.n9 stage1.n2 741
R362 stage1.n6 stage1.n2 741
R363 stage1.n7 stage1.n6 741
R364 stage1.n5 stage1.t0 323.575
R365 stage1.n9 stage1.n8 236.839
R366 stage1.n5 stage1.n4 151.427
R367 stage1.n3 stage1.n0 146.447
R368 stage1.n3 stage1.n1 146.447
R369 stage1.n10 stage1.n1 139.639
R370 stage1.n11 stage1.n0 133.804
R371 stage1 stage1.t1 69.0795
R372 stage1.n10 stage1.n9 46.2505
R373 stage1.n6 stage1.n3 46.2505
R374 stage1.n6 stage1.n5 46.2505
R375 stage1.n7 stage1.n1 46.2505
R376 stage1.n2 stage1.n0 46.2505
R377 stage1.t0 stage1.n2 46.2505
R378 stage1.n8 stage1.n7 29.6199
R379 stage1.n8 stage1.t0 14.7834
R380 stage1.n12 stage1.n11 5.56832
R381 stage1.n11 stage1.n10 3.2005
R382 stage1 stage1.n12 3.063
R383 stage1.n12 stage1.t2 1.84196
C0 VPWR vout 0.118949f
C1 clk ena 0.034743f
C2 m2_3648_12070# m2_2864_8934# 0.135204f
C3 ui_in[3] ui_in[2] 0.031023f
C4 stage3 stage2 1.1489f
C5 uio_in[4] uio_in[3] 0.031023f
C6 VPWR uio_in[3] 1.03e-19
C7 m2_3648_12070# m2_3592_15598# 0.104769f
C8 VPWR ui_in[1] 1.03e-19
C9 ui_in[5] VPWR 1.03e-19
C10 m2_3592_4230# m2_1800_4342# 0.559432f
C11 VPWR ui_in[0] 1.03e-19
C12 ui_in[0] ui_in[1] 0.031023f
C13 VPWR ui_in[4] 1.03e-19
C14 clk clka 0.366934f
C15 uio_in[1] uio_in[2] 0.031023f
C16 VPWR ui_in[7] 1.03e-19
C17 ui_in[5] ui_in[4] 0.031023f
C18 stage3 clkb 0.080496f
C19 m2_2472_13022# m2_3648_12070# 0.105624f
C20 VPWR clkb 1.72951f
C21 clkb stage2 57.2718f
C22 uio_in[7] uio_in[6] 0.031023f
C23 stage1 VPWR 0.51574f
C24 stage1 stage2 1.20983f
C25 VPWR ui_in[2] 1.03e-19
C26 rst_n clka 3.03e-19
C27 ui_in[2] ui_in[1] 0.031023f
C28 m2_2584_17838# m2_3592_15598# 0.151985f
C29 m2_1800_4342# m2_2864_8934# 0.00172f
C30 m2_3592_27358# m2_2584_29654# 0.091013f
C31 m2_3592_35982# m2_3592_39062# 0.162853f
C32 stage3 clka 57.1062f
C33 clka vout 0.021853f
C34 stage1 clkb 0.165327f
C35 VPWR clka 4.89721f
C36 uio_in[1] VPWR 1.03e-19
C37 stage2 clka 0.216306f
C38 VPWR uio_in[0] 1.03e-19
C39 rst_n clk 0.031944f
C40 ua[0] vout 12.5848f
C41 m2_1800_4342# ua[6] 0.004395f
C42 VPWR ua[0] 0.268291f
C43 VPWR ui_in[6] 1.03e-19
C44 uio_in[4] uio_in[5] 0.031023f
C45 ui_in[5] ui_in[6] 0.031023f
C46 ui_in[7] uio_in[0] 0.031023f
C47 VPWR uio_in[2] 1.03e-19
C48 VPWR clk 0.404729f
C49 uio_in[2] uio_in[3] 0.031023f
C50 clkb clka 2.835f
C51 ui_in[7] ui_in[6] 0.031023f
C52 stage1 clka 57.232803f
C53 clk ui_in[1] 2.07e-20
C54 m2_2808_33406# m2_2584_29654# 0.041637f
C55 VPWR ui_in[3] 1.03e-19
C56 clk ui_in[0] 9.82e-20
C57 uio_in[6] uio_in[5] 0.031023f
C58 m2_3592_27358# m2_2864_23326# 0.138713f
C59 m2_3592_42086# m2_3592_39062# 0.130452f
C60 ua[1] ua[0] 0.001614f
C61 ui_in[3] ui_in[4] 0.031023f
C62 VPWR rst_n 1.03e-19
C63 m2_2808_33406# m2_3592_35982# 0.0711f
C64 rst_n ui_in[0] 0.031023f
C65 m2_2472_13022# m2_2864_8934# 0.017782f
C66 stage3 vout 0.416737f
C67 uio_in[1] uio_in[0] 0.031023f
C68 ua[1] VGND 0.145965f
C69 ua[2] VGND 0.148302f
C70 ua[3] VGND 0.148302f
C71 ua[4] VGND 0.148302f
C72 ua[5] VGND 0.148302f
C73 ua[6] VGND 0.142703f
C74 ua[7] VGND 0.146962f
C75 ena VGND 0.075936f
C76 rst_n VGND 0.04853f
C77 ui_in[0] VGND 0.048746f
C78 ui_in[1] VGND 0.048746f
C79 ui_in[2] VGND 0.048746f
C80 ui_in[3] VGND 0.048746f
C81 ui_in[4] VGND 0.048746f
C82 ui_in[5] VGND 0.048746f
C83 ui_in[6] VGND 0.048746f
C84 ui_in[7] VGND 0.048746f
C85 uio_in[0] VGND 0.048746f
C86 uio_in[1] VGND 0.048746f
C87 uio_in[2] VGND 0.048746f
C88 uio_in[3] VGND 0.048746f
C89 uio_in[4] VGND 0.048746f
C90 uio_in[5] VGND 0.048746f
C91 uio_in[6] VGND 0.048746f
C92 uio_in[7] VGND 0.079769f
C93 clk VGND 1.75558f
C94 ua[0] VGND 45.063232f
C95 VPWR VGND 25.824959f
C96 m2_3592_4230# VGND 2.41736f $ **FLOATING
C97 m2_1800_4342# VGND 11.662f $ **FLOATING
C98 m2_2864_8934# VGND 5.1283f $ **FLOATING
C99 m2_3648_12070# VGND 3.18023f $ **FLOATING
C100 m2_2472_13022# VGND 0.831538f $ **FLOATING
C101 m2_3592_15598# VGND 5.94344f $ **FLOATING
C102 m2_2584_17838# VGND 4.71527f $ **FLOATING
C103 m2_2864_23326# VGND 4.89346f $ **FLOATING
C104 m2_3592_27358# VGND 4.41841f $ **FLOATING
C105 m2_2584_29654# VGND 4.17312f $ **FLOATING
C106 m2_2808_33406# VGND 4.18017f $ **FLOATING
C107 m2_3592_35982# VGND 4.2612f $ **FLOATING
C108 m2_3592_39062# VGND 5.95916f $ **FLOATING
C109 m2_3592_42086# VGND 4.32567f $ **FLOATING
C110 clkb VGND 17.0008f
C111 clka VGND 32.465546f
C112 vout VGND 0.123462p
C113 stage3 VGND 6.026126f
C114 stage2 VGND 6.755722f
C115 stage1 VGND 7.464655f
C116 stage1.t2 VGND 54.924603f
C117 stage1.n0 VGND 0.014847f
C118 stage1.n1 VGND 0.015108f
C119 stage1.n2 VGND 0.026122f
C120 stage1.t0 VGND 0.151293f
C121 stage1.n3 VGND 0.015426f
C122 stage1.n4 VGND 0.031578f
C123 stage1.n5 VGND 0.099057f
C124 stage1.n6 VGND 0.026411f
C125 stage1.n7 VGND 0.026122f
C126 stage1.n9 VGND 0.140709f
C127 stage1.n10 VGND 0.009264f
C128 stage1.n11 VGND 0.024349f
C129 stage1.n12 VGND 0.705173f
C130 stage1.t1 VGND 0.052067f
C131 VPWR.t1 VGND 0.004897f
C132 VPWR.n0 VGND 0.01181f
C133 VPWR.t2 VGND 0.004894f
C134 VPWR.n1 VGND 0.005048f
C135 VPWR.n2 VGND 0.005251f
C136 VPWR.n3 VGND 0.005251f
C137 VPWR.n4 VGND 0.005251f
C138 VPWR.t0 VGND 0.084375f
C139 VPWR.n5 VGND 0.005251f
C140 VPWR.n6 VGND 0.005251f
C141 VPWR.n7 VGND 0.002595f
C142 VPWR.n8 VGND 0.004931f
C143 VPWR.n9 VGND 0.00517f
C144 VPWR.n10 VGND 0.00517f
C145 VPWR.n11 VGND 0.065974f
C146 VPWR.n12 VGND 0.00517f
C147 VPWR.n13 VGND 0.00517f
C148 VPWR.n14 VGND 0.005251f
C149 VPWR.n15 VGND 0.002895f
C150 VPWR.n16 VGND 0.00517f
C151 VPWR.n17 VGND 0.065974f
C152 VPWR.n18 VGND 0.00517f
C153 VPWR.n19 VGND 0.002782f
C154 VPWR.n20 VGND 0.002591f
C155 VPWR.n21 VGND 0.007181f
C156 VPWR.n22 VGND 0.020781f
C157 VPWR.t3 VGND 0.021432f
C158 VPWR.n23 VGND 2.43955f
C159 stage3.t2 VGND 0.051318f
C160 stage3.t1 VGND 55.3166f
C161 stage3.n0 VGND 0.015024f
C162 stage3.n1 VGND 0.01533f
C163 stage3.n2 VGND 0.026303f
C164 stage3.t0 VGND 0.152337f
C165 stage3.n3 VGND 0.015532f
C166 stage3.n4 VGND 0.031796f
C167 stage3.n5 VGND 0.09974f
C168 stage3.n6 VGND 0.026593f
C169 stage3.n7 VGND 0.026303f
C170 stage3.n9 VGND 0.14168f
C171 stage3.n10 VGND 0.008747f
C172 stage3.n11 VGND 0.046769f
C173 stage3.n12 VGND 0.429482f
C174 stage3.n13 VGND 0.266759f
C175 vout.t2 VGND 8.12866f
C176 vout.n0 VGND 0.003396f
C177 vout.n1 VGND 0.003427f
C178 vout.n2 VGND 0.005837f
C179 vout.n3 VGND 0.005837f
C180 vout.n4 VGND 0.003447f
C181 vout.n5 VGND 0.031442f
C182 vout.t3 VGND 0.033807f
C183 vout.n7 VGND 0.007056f
C184 vout.n8 VGND 0.022135f
C185 vout.n9 VGND 0.005902f
C186 vout.n10 VGND 0.002228f
C187 vout.n11 VGND 0.080331f
C188 vout.n12 VGND 0.912319f
C189 vout.t1 VGND 0.001136f
C190 vout.n13 VGND 0.036828f
C191 vout.n14 VGND 0.037218f
C192 vout.n16 VGND 0.063332f
C193 vout.n17 VGND 0.037476f
C194 vout.n18 VGND 0.429581f
C195 vout.t0 VGND 0.70815f
C196 vout.n20 VGND 0.063332f
C197 vout.n21 VGND 0.429581f
C198 vout.n22 VGND 0.019117f
C199 vout.n23 VGND 0.018772f
C200 vout.n24 VGND 0.236039f
C201 ua[0].t1 VGND 0.005268f
C202 ua[0].t0 VGND 2.96209f
C203 ua[0].n0 VGND 0.263857f
C204 ua[0].t3 VGND 0.005265f
C205 ua[0].n1 VGND 0.025355f
C206 ua[0].n2 VGND 0.013735f
C207 ua[0].n3 VGND 0.173955f
C208 ua[0].n5 VGND 1.99399f
C209 ua[0].n6 VGND 0.087333f
C210 ua[0].n7 VGND 0.166073f
C211 ua[0].n8 VGND 0.293969f
C212 ua[0].t2 VGND 3.28704f
C213 ua[0].n10 VGND 1.99399f
C214 ua[0].n11 VGND 0.293969f
C215 ua[0].n12 VGND 0.166073f
C216 ua[0].n13 VGND 0.086792f
C217 ua[0].n14 VGND 0.014191f
C218 ua[0].n15 VGND 0.086114f
C219 clkb.t0 VGND 58.603302f
C220 clkb.t2 VGND 0.020864f
C221 clkb.t1 VGND 0.032902f
C222 stage2.t1 VGND 55.0583f
C223 stage2.n0 VGND 0.014797f
C224 stage2.n1 VGND 0.014928f
C225 stage2.n2 VGND 0.026188f
C226 stage2.t0 VGND 0.151672f
C227 stage2.n3 VGND 0.015465f
C228 stage2.n4 VGND 0.031658f
C229 stage2.n5 VGND 0.099305f
C230 stage2.n6 VGND 0.026477f
C231 stage2.n7 VGND 0.026188f
C232 stage2.n9 VGND 0.141061f
C233 stage2.n10 VGND 0.010925f
C234 stage2.n11 VGND 0.02724f
C235 stage2.n12 VGND 0.690044f
C236 stage2.t2 VGND 0.052779f
C237 clka.t2 VGND 0.080535f
C238 clka.t1 VGND 59.9508f
C239 clka.t0 VGND 58.621803f
C240 clka.n0 VGND 2.92909f
.ends

