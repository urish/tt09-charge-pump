* Dickson Charge Pump Teshbench
* Run with `make sim_nand`

.include "pdk_lib.spice"

* Power supply
V1 VGND 0 0
V2 VDPWR VGND 1.8
V3 VAPWR VGND 3.3
* Clock
V4 clk VGND PULSE(0 1.8 0 0 0 250n 500n)

.include "tt_um_urish_charge_pump.spice"

x1 clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
+ VGND VGND VGND VGND VGND VGND VGND VGND
+ VGND VGND VGND VGND VGND VGND VGND VGND
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VAPWR VGND VDPWR
+ tt_um_urish_charge_pump

.tran 10n 30u

.control
run
plot "ua[0]" x1.vout clk x1.stage1.t0 x1.stage2.t0 x1.stage3.t0
.endc
.end

.end
