magic
tech sky130A
magscale 1 2
timestamp 1725613538
<< error_s >>
rect 29099 44801 29100 44860
rect 799 44741 859 44801
rect 29100 44699 29101 44800
<< dnwell >>
rect 19800 40800 22260 43080
rect 19800 35460 22260 37740
rect 19800 30000 22260 32280
rect 19800 26400 22260 28680
<< nwell >>
rect 19720 42874 22340 43160
rect 19720 41006 20006 42874
rect 22054 41006 22340 42874
rect 19720 40720 22340 41006
rect 19720 37534 22340 37820
rect 19720 35666 20006 37534
rect 22054 35666 22340 37534
rect 19720 35380 22340 35666
rect 19720 32074 22340 32360
rect 19720 30206 20006 32074
rect 22054 30206 22340 32074
rect 19720 29920 22340 30206
rect 19720 28474 22340 28760
rect 19720 26606 20006 28474
rect 22054 26606 22340 28474
rect 19720 26320 22340 26606
<< nsubdiff >>
rect 19757 43103 22303 43123
rect 19757 43069 19837 43103
rect 22223 43069 22303 43103
rect 19757 43049 22303 43069
rect 19757 43043 19831 43049
rect 19757 40837 19777 43043
rect 19811 40837 19831 43043
rect 19757 40831 19831 40837
rect 22229 43043 22303 43049
rect 22229 40837 22249 43043
rect 22283 40837 22303 43043
rect 22229 40831 22303 40837
rect 19757 40811 22303 40831
rect 19757 40777 19837 40811
rect 22223 40777 22303 40811
rect 19757 40757 22303 40777
rect 19757 37763 22303 37783
rect 19757 37729 19837 37763
rect 22223 37729 22303 37763
rect 19757 37709 22303 37729
rect 19757 37703 19831 37709
rect 19757 35497 19777 37703
rect 19811 35497 19831 37703
rect 19757 35491 19831 35497
rect 22229 37703 22303 37709
rect 22229 35497 22249 37703
rect 22283 35497 22303 37703
rect 22229 35491 22303 35497
rect 19757 35471 22303 35491
rect 19757 35437 19837 35471
rect 22223 35437 22303 35471
rect 19757 35417 22303 35437
rect 19757 32303 22303 32323
rect 19757 32269 19837 32303
rect 22223 32269 22303 32303
rect 19757 32249 22303 32269
rect 19757 32243 19831 32249
rect 19757 30037 19777 32243
rect 19811 30037 19831 32243
rect 19757 30031 19831 30037
rect 22229 32243 22303 32249
rect 22229 30037 22249 32243
rect 22283 30037 22303 32243
rect 22229 30031 22303 30037
rect 19757 30011 22303 30031
rect 19757 29977 19837 30011
rect 22223 29977 22303 30011
rect 19757 29957 22303 29977
rect 19757 28703 22303 28723
rect 19757 28669 19837 28703
rect 22223 28669 22303 28703
rect 19757 28649 22303 28669
rect 19757 28643 19831 28649
rect 19757 26437 19777 28643
rect 19811 26437 19831 28643
rect 19757 26431 19831 26437
rect 22229 28643 22303 28649
rect 22229 26437 22249 28643
rect 22283 26437 22303 28643
rect 22229 26431 22303 26437
rect 19757 26411 22303 26431
rect 19757 26377 19837 26411
rect 22223 26377 22303 26411
rect 19757 26357 22303 26377
<< nsubdiffcont >>
rect 19837 43069 22223 43103
rect 19777 40837 19811 43043
rect 22249 40837 22283 43043
rect 19837 40777 22223 40811
rect 19837 37729 22223 37763
rect 19777 35497 19811 37703
rect 22249 35497 22283 37703
rect 19837 35437 22223 35471
rect 19837 32269 22223 32303
rect 19777 30037 19811 32243
rect 22249 30037 22283 32243
rect 19837 29977 22223 30011
rect 19837 28669 22223 28703
rect 19777 26437 19811 28643
rect 22249 26437 22283 28643
rect 19837 26377 22223 26411
<< locali >>
rect 31012 43728 31070 43762
rect 19777 43069 19837 43103
rect 22223 43069 22283 43103
rect 19777 43043 19811 43069
rect 22249 43043 22283 43069
rect 19777 40811 19811 40837
rect 22249 40811 22283 40837
rect 19777 40777 19837 40811
rect 22223 40777 22283 40811
rect 19777 37729 19837 37763
rect 22223 37729 22283 37763
rect 19777 37703 19811 37729
rect 22249 37703 22283 37729
rect 19777 35471 19811 35497
rect 22249 35471 22283 35497
rect 19777 35437 19837 35471
rect 22223 35437 22283 35471
rect 19777 32269 19837 32303
rect 22223 32269 22283 32303
rect 19777 32243 19811 32269
rect 22249 32243 22283 32269
rect 19777 30011 19811 30037
rect 22249 30011 22283 30037
rect 19777 29977 19837 30011
rect 22223 29977 22283 30011
rect 19777 28669 19837 28703
rect 22223 28669 22283 28703
rect 19777 28643 19811 28669
rect 22249 28643 22283 28669
rect 19777 26411 19811 26437
rect 22249 26411 22283 26437
rect 19777 26377 19837 26411
rect 22223 26377 22283 26411
<< viali >>
rect 30512 44468 30570 44502
rect 31012 44466 31070 44500
rect 30336 44280 30370 44340
rect 31212 44302 31246 44356
rect 30336 43620 30370 43680
rect 31212 43542 31246 43596
rect 20040 43103 20280 43140
rect 20040 43080 20280 43103
rect 20160 42780 20280 42840
rect 20160 37763 20340 37800
rect 20160 37729 20340 37763
rect 20160 37680 20340 37729
rect 20160 37440 20340 37500
rect 20160 31980 20340 32040
rect 21780 28703 21960 28740
rect 21780 28669 21960 28703
rect 21780 28620 21960 28669
rect 21780 28380 21900 28440
rect 23276 2902 23312 2948
rect 31490 1966 31530 2000
rect 31490 1478 31530 1512
<< metal1 >>
rect 30500 44502 30760 44520
rect 30500 44468 30512 44502
rect 30570 44468 30760 44502
rect 30500 44460 30760 44468
rect 30820 44506 31080 44520
rect 30820 44500 31082 44506
rect 30820 44466 31012 44500
rect 31070 44466 31082 44500
rect 30820 44460 31082 44466
rect 31200 44360 31260 44520
rect 30330 44340 30376 44352
rect 29150 44280 29160 44340
rect 29340 44280 30336 44340
rect 30370 44280 30480 44340
rect 30580 44300 31000 44360
rect 31100 44356 31260 44360
rect 31100 44302 31212 44356
rect 31246 44302 31260 44356
rect 31100 44300 31260 44302
rect 30330 44268 30376 44280
rect 30760 43980 30820 44300
rect 30750 43920 30760 43980
rect 30820 43920 30830 43980
rect 30760 43780 30820 43920
rect 30480 43720 31100 43780
rect 30330 43680 30376 43692
rect 29150 43620 29160 43680
rect 29340 43620 30336 43680
rect 30370 43620 30480 43680
rect 30330 43608 30376 43620
rect 31200 43600 31260 44300
rect 30600 43540 30980 43600
rect 31100 43596 31260 43600
rect 31100 43542 31212 43596
rect 31246 43542 31260 43596
rect 31100 43540 31260 43542
rect 20030 43260 20040 43440
rect 20280 43260 20290 43440
rect 20040 43146 20280 43260
rect 20028 43140 20292 43146
rect 30680 43140 30740 43540
rect 31200 43400 31260 43540
rect 31190 43280 31200 43400
rect 31260 43280 31270 43400
rect 20028 43080 20040 43140
rect 20280 43080 20292 43140
rect 20028 43074 20292 43080
rect 20040 42846 20280 43074
rect 30650 42960 30660 43140
rect 30780 42960 30790 43140
rect 20040 42840 20292 42846
rect 20040 42780 20160 42840
rect 20280 42780 20292 42840
rect 20040 42774 20292 42780
rect 20040 42540 20280 42774
rect 21840 42120 22320 42300
rect 22500 42120 22510 42300
rect 20150 37860 20160 38040
rect 20340 37860 20350 38040
rect 20160 37806 20340 37860
rect 20148 37800 20352 37806
rect 20148 37680 20160 37800
rect 20340 37680 20352 37800
rect 20148 37674 20352 37680
rect 20160 37506 20340 37674
rect 20148 37500 20352 37506
rect 20148 37440 20160 37500
rect 20340 37440 20352 37500
rect 20148 37434 20352 37440
rect 20160 37140 20340 37434
rect 21840 36480 22320 36660
rect 22500 36480 22510 36660
rect 20150 32400 20160 32580
rect 20340 32400 20350 32580
rect 20160 32046 20340 32400
rect 20148 32040 20352 32046
rect 20148 31980 20160 32040
rect 20340 31980 20352 32040
rect 20148 31974 20352 31980
rect 20160 31680 20340 31974
rect 21840 31242 22514 31260
rect 21840 31096 22362 31242
rect 22498 31096 22514 31242
rect 21840 31080 22514 31096
rect 21770 28800 21780 28980
rect 21960 28800 21970 28980
rect 21780 28746 21960 28800
rect 21768 28740 21972 28746
rect 21768 28620 21780 28740
rect 21960 28620 21972 28740
rect 21768 28614 21972 28620
rect 21780 28446 21960 28614
rect 21768 28440 21960 28446
rect 21768 28380 21780 28440
rect 21900 28380 21960 28440
rect 21768 28374 21960 28380
rect 19380 28140 20220 28200
rect 19370 27900 19380 28140
rect 19620 27900 20220 28140
rect 21780 28080 21960 28374
rect 19380 27660 20220 27900
rect 19370 27420 19380 27660
rect 19620 27420 20220 27660
rect 19380 27180 20220 27420
rect 19370 26940 19380 27180
rect 19620 26940 20220 27180
rect 19380 26880 20220 26940
rect 23060 2898 23070 2960
rect 23126 2948 23136 2960
rect 23270 2948 23318 2960
rect 23126 2902 23276 2948
rect 23312 2902 23429 2948
rect 23126 2898 23136 2902
rect 23270 2890 23318 2902
rect 23383 2793 23429 2902
rect 31490 2752 31530 2902
rect 31442 2706 31530 2752
rect 31490 2392 31530 2706
rect 31460 2246 31470 2392
rect 31538 2246 31548 2392
rect 31490 2006 31530 2246
rect 31478 2000 31542 2006
rect 31478 1966 31490 2000
rect 31530 1966 31542 2000
rect 31478 1960 31542 1966
rect 23394 1132 23496 1864
rect 31490 1518 31530 1960
rect 31478 1512 31542 1518
rect 31478 1478 31490 1512
rect 31530 1478 31542 1512
rect 31478 1472 31542 1478
rect 23394 1032 23404 1132
rect 23488 1032 23498 1132
rect 23394 1020 23496 1032
<< via1 >>
rect 30760 44460 30820 44520
rect 29160 44280 29340 44340
rect 30760 43920 30820 43980
rect 29160 43620 29340 43680
rect 20040 43260 20280 43440
rect 31200 43280 31260 43400
rect 30660 42960 30780 43140
rect 22320 42120 22500 42300
rect 20160 37860 20340 38040
rect 22320 36480 22500 36660
rect 20160 32400 20340 32580
rect 22362 31096 22498 31242
rect 21780 28800 21960 28980
rect 19380 27900 19620 28140
rect 19380 27420 19620 27660
rect 19380 26940 19620 27180
rect 23070 2898 23126 2960
rect 31470 2246 31538 2392
rect 23404 1032 23488 1132
<< metal2 >>
rect 28750 45042 28850 45052
rect 28750 44932 28850 44942
rect 28770 44882 28830 44932
rect 28770 44822 30820 44882
rect 30760 44520 30820 44822
rect 30760 44450 30820 44460
rect 29160 44340 29340 44350
rect 29160 44270 29340 44280
rect 27900 43980 28020 43990
rect 30760 43980 30820 43990
rect 28020 43920 30760 43980
rect 30820 43920 30840 43980
rect 28020 43860 30840 43920
rect 27900 43850 28020 43860
rect 29160 43680 29340 43690
rect 29160 43610 29340 43620
rect 20040 43440 20280 43450
rect 20040 43250 20280 43260
rect 22320 42300 22500 42310
rect 20160 38040 20340 38050
rect 22320 38040 22500 42120
rect 20340 37860 22500 38040
rect 20160 37850 20340 37860
rect 22320 37800 22500 37860
rect 22320 36660 22500 36670
rect 20160 32580 20340 32590
rect 22320 32580 22500 36480
rect 20340 32400 22500 32580
rect 20160 32390 20340 32400
rect 29580 32040 29700 43860
rect 31200 43400 31260 43410
rect 31200 43270 31260 43280
rect 30660 43140 30780 43150
rect 30660 42950 30780 42960
rect 29580 31910 29700 31920
rect 22336 31242 22516 31256
rect 22336 31096 22362 31242
rect 22498 31096 22516 31242
rect 21780 28980 21960 28990
rect 22336 28980 22516 31096
rect 21960 28800 22516 28980
rect 21780 28790 21960 28800
rect 19380 28140 19620 28150
rect 19380 27890 19620 27900
rect 19380 27660 19620 27670
rect 19380 27410 19620 27420
rect 19380 27180 19620 27190
rect 19380 26930 19620 26940
rect 23070 2960 23126 2970
rect 23070 2888 23126 2898
rect 31470 2392 31538 2402
rect 31470 2236 31538 2246
rect 9900 1140 10020 1150
rect 23404 1140 23488 1142
rect 10020 1132 23494 1140
rect 10020 1032 23404 1132
rect 23488 1032 23494 1132
rect 10020 1020 23494 1032
rect 9900 1010 10020 1020
<< via2 >>
rect 28750 44942 28850 45042
rect 29160 44280 29340 44340
rect 27900 43860 28020 43980
rect 29160 43620 29340 43680
rect 20040 43260 20280 43440
rect 22320 42120 22500 42300
rect 22320 36480 22500 36660
rect 31200 43280 31260 43400
rect 30660 42960 30780 43140
rect 29580 31920 29700 32040
rect 22362 31096 22498 31242
rect 19380 27900 19620 28140
rect 19380 27420 19620 27660
rect 19380 26940 19620 27180
rect 23070 2898 23126 2960
rect 31470 2246 31538 2392
rect 9900 1020 10020 1140
<< metal3 >>
rect 28740 45042 28860 45047
rect 28740 44942 28750 45042
rect 28850 44942 28860 45042
rect 28740 44937 28860 44942
rect 29090 44500 29100 44800
rect 29400 44500 29410 44800
rect 29100 44340 29400 44500
rect 29100 44280 29160 44340
rect 29340 44280 29400 44340
rect 27890 43980 28030 43985
rect 27890 43860 27900 43980
rect 28020 43860 28030 43980
rect 27890 43855 28030 43860
rect 29100 43680 29400 44280
rect 20130 43500 28640 43680
rect 29100 43620 29160 43680
rect 29340 43620 29400 43680
rect 29100 43600 29400 43620
rect 20130 43445 20310 43500
rect 20030 43440 20310 43445
rect 28460 43440 28640 43500
rect 20030 43260 20040 43440
rect 20280 43260 20310 43440
rect 28432 43260 28440 43440
rect 28740 43400 28750 43440
rect 31190 43400 31270 43405
rect 28740 43280 31200 43400
rect 31260 43280 31270 43400
rect 28740 43260 28750 43280
rect 31190 43275 31270 43280
rect 20030 43255 20310 43260
rect 28460 43246 28640 43260
rect 30650 43140 30790 43145
rect 30650 42960 30660 43140
rect 30780 42960 30790 43140
rect 30650 42955 30790 42960
rect 22310 42300 22510 42305
rect 22310 42120 22320 42300
rect 22500 42120 22510 42300
rect 22310 42115 22510 42120
rect 30660 37440 30780 42955
rect 28070 37320 28080 37440
rect 28260 37320 30780 37440
rect 22310 36660 22510 36665
rect 22310 36480 22320 36660
rect 22500 36480 22510 36660
rect 22310 36475 22510 36480
rect 29570 32040 29710 32045
rect 28070 31920 28080 32040
rect 28260 31920 29580 32040
rect 29700 31920 29710 32040
rect 29570 31915 29710 31920
rect 22352 31242 22508 31247
rect 22352 31096 22362 31242
rect 22498 31096 22508 31242
rect 22352 31091 22508 31096
rect 19380 28145 19620 28200
rect 19370 28140 19630 28145
rect 19370 27900 19380 28140
rect 19620 27900 19630 28140
rect 19370 27895 19630 27900
rect 19380 27665 19620 27895
rect 19370 27660 19630 27665
rect 19370 27420 19380 27660
rect 19620 27420 19630 27660
rect 19370 27415 19630 27420
rect 19380 27185 19620 27415
rect 19370 27180 19630 27185
rect 19370 26940 19380 27180
rect 19620 26940 19630 27180
rect 19370 26935 19630 26940
rect 19380 3136 19620 26935
rect 19380 2965 23130 3136
rect 19380 2960 23136 2965
rect 19380 2898 23070 2960
rect 23126 2898 23136 2960
rect 19380 2896 23136 2898
rect 23060 2893 23136 2896
rect 31460 2392 31548 2397
rect 31460 2246 31470 2392
rect 31538 2246 31548 2392
rect 31460 2241 31548 2246
rect 9890 1140 10030 1145
rect 9890 1020 9900 1140
rect 10020 1020 10030 1140
rect 9890 1015 10030 1020
<< via3 >>
rect 28750 44942 28850 45042
rect 29100 44500 29400 44800
rect 27900 43860 28020 43980
rect 28440 43260 28740 43440
rect 22320 42120 22500 42300
rect 28080 37320 28260 37440
rect 22320 36480 22500 36660
rect 28080 31920 28260 32040
rect 22362 31096 22498 31242
rect 19380 27900 19620 28140
rect 19380 27420 19620 27660
rect 19380 26940 19620 27180
rect 31470 2246 31538 2392
rect 9900 1020 10020 1140
<< metal4 >>
rect 799 44741 800 44801
rect 6134 44700 6194 45152
rect 6686 44700 6746 45152
rect 7238 44700 7298 45152
rect 7790 44700 7850 45152
rect 8342 44700 8402 45152
rect 8894 44700 8954 45152
rect 9446 44700 9506 45152
rect 9998 44700 10058 45152
rect 10550 44700 10610 45152
rect 11102 44700 11162 45152
rect 11654 44700 11714 45152
rect 12206 44700 12266 45152
rect 12758 44700 12818 45152
rect 13310 44700 13370 45152
rect 13862 44700 13922 45152
rect 14414 44700 14474 45152
rect 14966 44700 15026 45152
rect 15518 44700 15578 45152
rect 16070 44700 16130 45152
rect 16622 44700 16682 45152
rect 17174 44700 17234 45152
rect 17726 44700 17786 45152
rect 18278 44700 18338 45152
rect 18830 44700 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 45043 28826 45152
rect 28749 45042 28851 45043
rect 28749 44942 28750 45042
rect 28850 44942 28851 45042
rect 29318 44952 29378 45152
rect 28749 44941 28851 44942
rect 29099 44800 29401 44801
rect 6126 44500 29100 44700
rect 29400 44500 29401 44800
rect 9800 27840 10100 44500
rect 29099 44499 29401 44500
rect 27899 43980 28021 43981
rect 27899 43860 27900 43980
rect 28020 43860 28021 43980
rect 27899 43859 28021 43860
rect 27900 43020 28020 43859
rect 28440 43441 28740 44152
rect 28439 43440 28741 43441
rect 28439 43260 28440 43440
rect 28740 43260 28741 43440
rect 28439 43259 28741 43260
rect 22319 42300 22501 42301
rect 22319 42120 22320 42300
rect 22500 42120 22920 42300
rect 22319 42119 22501 42120
rect 27900 37440 28320 37620
rect 27900 37320 28080 37440
rect 28260 37320 28320 37440
rect 27900 37200 28320 37320
rect 22319 36660 22501 36661
rect 22319 36480 22320 36660
rect 22500 36480 22860 36660
rect 22319 36479 22501 36480
rect 27900 32040 28320 32160
rect 27900 31920 28080 32040
rect 28260 31920 28320 32040
rect 27900 31800 28320 31920
rect 22352 31242 22860 31260
rect 22352 31096 22362 31242
rect 22498 31096 22860 31242
rect 22352 31080 22860 31096
rect 19020 28141 19620 28200
rect 19020 28140 19621 28141
rect 19020 27900 19380 28140
rect 19620 27900 19621 28140
rect 19020 27899 19621 27900
rect 9800 25680 13080 27840
rect 19020 27661 19620 27899
rect 19020 27660 19621 27661
rect 19020 27420 19380 27660
rect 19620 27420 19621 27660
rect 19020 27419 19621 27420
rect 19020 27181 19620 27419
rect 19020 27180 19621 27181
rect 19020 26940 19380 27180
rect 19620 26940 19621 27180
rect 19020 26939 19621 26940
rect 19020 26880 19620 26939
rect 9800 1140 10100 25680
rect 9800 1020 9900 1140
rect 10020 1020 10100 1140
rect 9800 1000 10100 1020
rect 28440 1000 28740 43259
rect 31282 2392 31554 2408
rect 31282 2246 31470 2392
rect 31538 2246 31554 2392
rect 31282 2228 31554 2246
rect 31282 780 31462 2228
rect 30362 600 31462 780
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C1
timestamp 1711870259
transform 1 0 25350 0 1 40500
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C2
timestamp 1711870259
transform 1 0 25330 0 1 35060
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C3
timestamp 1711870259
transform 1 0 25330 0 1 29600
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_WMZ6NR  C4
timestamp 1711870259
transform 1 0 15990 0 1 26540
box -3150 -2600 3149 2600
use high_voltage_logo  high_voltage_logo_0
timestamp 1711967973
transform 0 -1 7568 1 0 1262
box 0 0 42336 5768
use sky130_fd_pr__pfet_01v8_BFP3TE  M1
timestamp 1711870259
transform 1 0 31041 0 1 44269
box -241 -369 241 369
use sky130_fd_pr__pfet_01v8_BFP3TE  M2
timestamp 1711870259
transform 1 0 31041 0 1 43531
box -241 -369 241 369
use sky130_fd_pr__nfet_01v8_DSY3K9  M3
timestamp 1711870259
transform -1 0 30541 0 1 44330
box -241 -310 241 310
use sky130_fd_pr__nfet_01v8_DSY3K9  M4
timestamp 1711870259
transform 1 0 30541 0 1 43592
box -241 -310 241 310
use sky130_fd_pr__nfet_01v8_lvt_WVNKYW  M5
timestamp 1711870259
transform 1 0 21036 0 1 41950
box -996 -910 996 910
use sky130_fd_pr__nfet_01v8_lvt_WVNKYW  M6
timestamp 1711870259
transform 1 0 21036 0 1 36610
box -996 -910 996 910
use sky130_fd_pr__nfet_01v8_lvt_WVNKYW  M7
timestamp 1711870259
transform 1 0 21036 0 1 31150
box -996 -910 996 910
use sky130_fd_pr__nfet_01v8_lvt_WVNKYW  M8
timestamp 1711870259
transform 1 0 21036 0 1 27550
box -996 -910 996 910
use sky130_fd_pr__pfet_g5v0d10v5_RSSSV2  M9
timestamp 1717238374
transform 1 0 27458 0 1 2835
box -4258 -339 4258 339
use sky130_fd_pr__pfet_g5v0d10v5_RSSSV2  M10
timestamp 1717238374
transform 1 0 27458 0 1 1739
box -4258 -339 4258 339
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal1 30760 43980 30820 44100 0 FreeSans 320 90 0 0 clka
flabel metal1 30680 42960 30740 43560 0 FreeSans 320 90 0 0 clkb
flabel metal2 22320 37800 22500 42120 0 FreeSans 1600 0 0 0 stage1
flabel metal2 22320 32400 22500 36480 0 FreeSans 1600 0 0 0 stage2
flabel metal3 19380 21660 19620 23880 0 FreeSans 1600 0 0 0 vout
flabel metal4 28440 1000 28740 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal2 22336 28800 22516 31080 0 FreeSans 1600 0 0 0 stage3
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
