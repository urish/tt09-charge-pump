magic
tech sky130A
magscale 1 2
timestamp 1725743120
<< viali >>
rect 27208 44280 27242 44340
rect 28268 44120 28304 44668
rect 27208 43620 27242 43680
rect 28268 43296 28304 43844
rect 18056 41780 18194 42604
rect 18708 42124 18756 42272
rect 18056 36156 18194 36980
rect 18714 36484 18776 36656
rect 18060 30744 18198 31568
rect 18716 31082 18756 31260
rect 18188 28248 18880 28342
rect 18296 27664 18356 28092
rect 28032 4170 28426 4214
rect 20250 3046 20530 3112
rect 28362 1966 28402 2000
rect 28362 1478 28402 1512
<< metal1 >>
rect 28154 44668 28316 44712
rect 27622 44626 27632 44636
rect 27405 44592 27632 44626
rect 27622 44584 27632 44592
rect 27692 44626 27702 44636
rect 27692 44592 28115 44626
rect 27692 44584 27702 44592
rect 27194 44340 27256 44360
rect 27298 44340 27358 44562
rect 27496 44414 28018 44474
rect 26022 44280 26032 44340
rect 26212 44280 27208 44340
rect 27242 44280 27358 44340
rect 27194 44250 27256 44280
rect 27632 43980 27692 44414
rect 28154 44120 28268 44668
rect 28304 44120 28316 44668
rect 27622 43920 27632 43980
rect 27692 43920 27702 43980
rect 27632 43832 27692 43920
rect 28154 43844 28316 44120
rect 27388 43772 28124 43832
rect 27202 43680 27248 43692
rect 26022 43620 26032 43680
rect 26212 43620 27208 43680
rect 27242 43620 27352 43680
rect 27202 43608 27248 43620
rect 27508 43566 28016 43600
rect 27504 43540 28016 43566
rect 27504 43524 27612 43540
rect 27552 43140 27612 43524
rect 28154 43392 28268 43844
rect 28154 43292 28222 43392
rect 28304 43296 28316 43844
rect 28278 43292 28316 43296
rect 28154 43284 28316 43292
rect 27522 42960 27532 43140
rect 27652 42960 27662 43140
rect 18050 42604 18200 42616
rect 18046 41780 18056 42604
rect 18194 41780 18204 42604
rect 18702 42274 18762 42284
rect 19038 42274 19192 42300
rect 18432 42104 18442 42274
rect 18612 42104 18622 42274
rect 18702 42272 19192 42274
rect 18702 42124 18708 42272
rect 18756 42124 19192 42272
rect 18702 42120 19192 42124
rect 19372 42120 19382 42300
rect 18702 42112 18762 42120
rect 18050 41768 18200 41780
rect 18050 36980 18200 36992
rect 18046 36156 18056 36980
rect 18194 36156 18204 36980
rect 18708 36660 18782 36668
rect 18708 36656 19192 36660
rect 18440 36476 18450 36656
rect 18630 36476 18640 36656
rect 18708 36484 18714 36656
rect 18776 36484 19192 36656
rect 18708 36480 19192 36484
rect 19372 36480 19382 36660
rect 18708 36472 18782 36480
rect 18050 36144 18200 36156
rect 18054 31568 18204 31580
rect 18050 30744 18060 31568
rect 18198 30744 18208 31568
rect 18710 31260 18762 31272
rect 18432 31074 18442 31246
rect 18614 31074 18624 31246
rect 18710 31082 18716 31260
rect 18756 31242 19386 31260
rect 18756 31096 19234 31242
rect 19370 31096 19386 31242
rect 18756 31082 19386 31096
rect 18710 31080 19386 31082
rect 18710 31070 18762 31080
rect 18054 30732 18204 30744
rect 18016 28354 19000 28356
rect 18014 28226 18024 28354
rect 18208 28342 19000 28354
rect 18880 28248 19000 28342
rect 18208 28226 19000 28248
rect 18016 28212 19000 28226
rect 16252 28146 17092 28200
rect 16252 28140 18368 28146
rect 16242 27900 16252 28140
rect 16492 28092 18368 28140
rect 16492 27900 18296 28092
rect 16252 27664 18296 27900
rect 18356 27664 18368 28092
rect 18430 27786 18440 27966
rect 18620 27786 18630 27966
rect 16252 27660 18368 27664
rect 16242 27420 16252 27660
rect 16492 27610 18368 27660
rect 16492 27420 17092 27610
rect 16252 27180 17092 27420
rect 16242 26940 16252 27180
rect 16492 26940 17092 27180
rect 16252 26880 17092 26940
rect 28314 4220 28324 4270
rect 28020 4214 28324 4220
rect 28516 4220 28526 4270
rect 28020 4170 28032 4214
rect 28020 4164 28324 4170
rect 28314 4152 28324 4164
rect 28516 4152 28528 4220
rect 20242 3118 20530 4078
rect 28356 3842 28528 4152
rect 20238 3112 20542 3118
rect 20238 3046 20250 3112
rect 20530 3046 20542 3112
rect 20238 3040 20542 3046
rect 20242 3010 20530 3040
rect 20242 2774 20292 3010
rect 28362 2752 28402 2902
rect 28314 2706 28402 2752
rect 28362 2392 28402 2706
rect 28332 2246 28342 2392
rect 28410 2246 28420 2392
rect 28362 2006 28402 2246
rect 28350 2000 28414 2006
rect 28350 1966 28362 2000
rect 28402 1966 28414 2000
rect 28350 1960 28414 1966
rect 20266 1132 20368 1864
rect 28362 1518 28402 1960
rect 28350 1512 28414 1518
rect 28350 1478 28362 1512
rect 28402 1478 28414 1512
rect 28350 1472 28414 1478
rect 20266 1032 20276 1132
rect 20360 1032 20370 1132
rect 20266 1020 20368 1032
<< via1 >>
rect 27632 44584 27692 44636
rect 26032 44280 26212 44340
rect 27632 43920 27692 43980
rect 26032 43620 26212 43680
rect 28222 43296 28268 43392
rect 28268 43296 28278 43392
rect 28222 43292 28278 43296
rect 27532 42960 27652 43140
rect 18056 41780 18194 42604
rect 18442 42104 18612 42274
rect 19192 42120 19372 42300
rect 18056 36156 18194 36980
rect 18450 36476 18630 36656
rect 19192 36480 19372 36660
rect 18060 30744 18198 31568
rect 18442 31074 18614 31246
rect 19234 31096 19370 31242
rect 18024 28342 18208 28354
rect 18024 28248 18188 28342
rect 18188 28248 18208 28342
rect 18024 28226 18208 28248
rect 16252 27900 16492 28140
rect 18440 27786 18620 27966
rect 16252 27420 16492 27660
rect 16252 26940 16492 27180
rect 28324 4214 28516 4270
rect 28324 4170 28426 4214
rect 28426 4170 28516 4214
rect 28324 4152 28516 4170
rect 28342 2246 28410 2392
rect 20276 1032 20360 1132
<< metal2 >>
rect 25622 45042 25722 45052
rect 25622 44932 25722 44942
rect 25642 44882 25702 44932
rect 25642 44822 27692 44882
rect 27632 44636 27692 44822
rect 27632 44574 27692 44584
rect 26032 44340 26212 44350
rect 26032 44270 26212 44280
rect 24772 43980 24892 43990
rect 27632 43980 27692 43990
rect 24892 43920 27632 43980
rect 27692 43920 27712 43980
rect 24892 43860 27712 43920
rect 24772 43850 24892 43860
rect 26032 43680 26212 43690
rect 26032 43610 26212 43620
rect 18056 42604 18194 42614
rect 19192 42300 19372 42310
rect 18442 42274 18612 42284
rect 18442 42094 18612 42104
rect 18056 41770 18194 41780
rect 19192 37344 19372 42120
rect 18434 37164 19372 37344
rect 18056 36980 18194 36990
rect 18434 36666 18614 37164
rect 18434 36656 18630 36666
rect 18434 36476 18450 36656
rect 18434 36474 18630 36476
rect 18450 36466 18630 36474
rect 19192 36660 19372 36670
rect 18056 36146 18194 36156
rect 19192 32132 19372 36480
rect 18434 31952 19372 32132
rect 26452 32040 26572 43860
rect 28222 43392 28278 43402
rect 28222 43282 28278 43292
rect 27532 43140 27652 43150
rect 27532 42950 27652 42960
rect 18060 31568 18198 31578
rect 18434 31246 18614 31952
rect 26452 31910 26572 31920
rect 18434 31074 18442 31246
rect 18434 31072 18614 31074
rect 18442 31064 18614 31072
rect 19208 31242 19388 31256
rect 19208 31096 19234 31242
rect 19370 31096 19388 31242
rect 18060 30734 18198 30744
rect 19208 28980 19388 31096
rect 18440 28800 19388 28980
rect 18024 28354 18208 28364
rect 18024 28216 18208 28226
rect 16252 28140 16492 28150
rect 16252 27890 16492 27900
rect 18440 27966 18620 28800
rect 18440 27776 18620 27786
rect 16252 27660 16492 27670
rect 16252 27410 16492 27420
rect 16252 27180 16492 27190
rect 16252 26930 16492 26940
rect 28324 4270 28516 4280
rect 28324 4142 28516 4152
rect 28342 2392 28410 2402
rect 28342 2236 28410 2246
rect 6772 1140 6892 1150
rect 20276 1140 20360 1142
rect 6892 1132 20366 1140
rect 6892 1032 20276 1132
rect 20360 1032 20366 1132
rect 6892 1020 20366 1032
rect 6772 1010 6892 1020
<< via2 >>
rect 25622 44942 25722 45042
rect 26032 44280 26212 44340
rect 24772 43860 24892 43980
rect 26032 43620 26212 43680
rect 18056 41780 18194 42604
rect 18442 42104 18612 42274
rect 19192 42120 19372 42300
rect 18056 36156 18194 36980
rect 19192 36480 19372 36660
rect 28222 43292 28278 43392
rect 27532 42960 27652 43140
rect 18060 30744 18198 31568
rect 26452 31920 26572 32040
rect 19234 31096 19370 31242
rect 18024 28226 18208 28354
rect 16252 27900 16492 28140
rect 16252 27420 16492 27660
rect 16252 26940 16492 27180
rect 28324 4152 28516 4270
rect 28342 2246 28410 2392
rect 6772 1020 6892 1140
<< metal3 >>
rect 25612 45042 25732 45047
rect 25612 44942 25622 45042
rect 25722 44942 25732 45042
rect 25612 44937 25732 44942
rect 25962 44500 25972 44700
rect 26272 44500 26282 44700
rect 25972 44340 26272 44500
rect 25972 44280 26032 44340
rect 26212 44280 26272 44340
rect 24762 43980 24902 43985
rect 24762 43860 24772 43980
rect 24892 43860 24902 43980
rect 24762 43855 24902 43860
rect 25972 43680 26272 44280
rect 18432 43500 25512 43680
rect 25972 43620 26032 43680
rect 26212 43620 26272 43680
rect 25972 43600 26272 43620
rect 18046 42604 18204 42609
rect 18046 41780 18056 42604
rect 18194 41780 18204 42604
rect 18432 42279 18612 43500
rect 25332 43440 25512 43500
rect 25304 43260 25312 43440
rect 25612 43400 25622 43440
rect 25612 43397 28286 43400
rect 25612 43392 28288 43397
rect 25612 43292 28222 43392
rect 28278 43292 28288 43392
rect 25612 43287 28288 43292
rect 25612 43280 28286 43287
rect 25612 43260 25622 43280
rect 25332 43246 25512 43260
rect 27522 43140 27662 43145
rect 27522 42960 27532 43140
rect 27652 42960 27662 43140
rect 27522 42955 27662 42960
rect 19182 42300 19382 42305
rect 18432 42274 18622 42279
rect 18432 42104 18442 42274
rect 18612 42104 18622 42274
rect 19182 42120 19192 42300
rect 19372 42120 19382 42300
rect 19182 42115 19382 42120
rect 18432 42099 18622 42104
rect 18432 42088 18612 42099
rect 18046 41775 18204 41780
rect 27532 37440 27652 42955
rect 24942 37320 24952 37440
rect 25132 37320 27652 37440
rect 18046 36980 18204 36985
rect 18046 36156 18056 36980
rect 18194 36156 18204 36980
rect 19182 36660 19382 36665
rect 19182 36480 19192 36660
rect 19372 36480 19382 36660
rect 19182 36475 19382 36480
rect 18046 36151 18204 36156
rect 26442 32040 26582 32045
rect 24942 31920 24952 32040
rect 25132 31920 26452 32040
rect 26572 31920 26582 32040
rect 26442 31915 26582 31920
rect 18050 31568 18208 31573
rect 18050 30744 18060 31568
rect 18198 30744 18208 31568
rect 19224 31242 19380 31247
rect 19224 31096 19234 31242
rect 19370 31096 19380 31242
rect 19224 31091 19380 31096
rect 18050 30739 18208 30744
rect 18014 28354 18218 28359
rect 18014 28226 18024 28354
rect 18208 28226 18218 28354
rect 18014 28221 18218 28226
rect 16252 28145 16492 28200
rect 16242 28140 16502 28145
rect 16242 27900 16252 28140
rect 16492 27900 16502 28140
rect 16242 27895 16502 27900
rect 16252 27665 16492 27895
rect 16242 27660 16502 27665
rect 16242 27420 16252 27660
rect 16492 27420 16502 27660
rect 16242 27415 16502 27420
rect 16252 27185 16492 27415
rect 16242 27180 16502 27185
rect 16242 26940 16252 27180
rect 16492 26940 16502 27180
rect 16242 26935 16502 26940
rect 16252 4994 16492 26935
rect 16252 4754 28538 4994
rect 28298 4270 28538 4754
rect 28298 4152 28324 4270
rect 28516 4152 28538 4270
rect 28298 4126 28538 4152
rect 28332 2392 28420 2397
rect 28332 2246 28342 2392
rect 28410 2246 28420 2392
rect 28332 2241 28420 2246
rect 6762 1140 6902 1145
rect 6762 1020 6772 1140
rect 6892 1020 6902 1140
rect 6762 1015 6902 1020
<< via3 >>
rect 25622 44942 25722 45042
rect 25972 44500 26272 44700
rect 24772 43860 24892 43980
rect 18056 41780 18194 42604
rect 25312 43260 25612 43440
rect 19192 42120 19372 42300
rect 24952 37320 25132 37440
rect 18056 36156 18194 36980
rect 19192 36480 19372 36660
rect 24952 31920 25132 32040
rect 18060 30744 18198 31568
rect 19234 31096 19370 31242
rect 18024 28226 18208 28354
rect 16252 27900 16492 28140
rect 16252 27420 16492 27660
rect 16252 26940 16492 27180
rect 28342 2246 28410 2392
rect 6772 1020 6892 1140
<< metal4 >>
rect 3006 44700 3066 45152
rect 3558 44700 3618 45152
rect 4110 44700 4170 45152
rect 4662 44700 4722 45152
rect 5214 44700 5274 45152
rect 5766 44700 5826 45152
rect 6318 44700 6378 45152
rect 6870 44700 6930 45152
rect 7422 44700 7482 45152
rect 7974 44700 8034 45152
rect 8526 44700 8586 45152
rect 9078 44700 9138 45152
rect 9630 44700 9690 45152
rect 10182 44700 10242 45152
rect 10734 44700 10794 45152
rect 11286 44700 11346 45152
rect 11838 44700 11898 45152
rect 12390 44700 12450 45152
rect 12942 44700 13002 45152
rect 13494 44700 13554 45152
rect 14046 44700 14106 45152
rect 14598 44700 14658 45152
rect 15150 44700 15210 45152
rect 15702 44700 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 45043 25698 45152
rect 25621 45042 25723 45043
rect 25621 44942 25622 45042
rect 25722 44942 25723 45042
rect 26190 44952 26250 45152
rect 25621 44941 25723 44942
rect 25971 44700 26273 44701
rect 2998 44500 25972 44700
rect 26272 44500 26273 44700
rect 6072 1000 6372 44152
rect 6672 27840 6972 44500
rect 18018 42604 18218 44500
rect 25971 44499 26273 44500
rect 24771 43980 24893 43981
rect 24771 43860 24772 43980
rect 24892 43860 24893 43980
rect 24771 43859 24893 43860
rect 24772 43020 24892 43859
rect 25312 43441 25612 44152
rect 25311 43440 25613 43441
rect 25311 43260 25312 43440
rect 25612 43260 25613 43440
rect 25311 43259 25613 43260
rect 18018 41780 18056 42604
rect 18194 41780 18218 42604
rect 19191 42300 19373 42301
rect 19191 42120 19192 42300
rect 19372 42120 19792 42300
rect 19191 42119 19373 42120
rect 18018 36980 18218 41780
rect 24772 37440 25192 37620
rect 24772 37320 24952 37440
rect 25132 37320 25192 37440
rect 24772 37200 25192 37320
rect 18018 36156 18056 36980
rect 18194 36156 18218 36980
rect 19191 36660 19373 36661
rect 19191 36480 19192 36660
rect 19372 36480 19732 36660
rect 19191 36479 19373 36480
rect 18018 31568 18218 36156
rect 24772 32040 25192 32160
rect 24772 31920 24952 32040
rect 25132 31920 25192 32040
rect 24772 31800 25192 31920
rect 18018 30744 18060 31568
rect 18198 30744 18218 31568
rect 19224 31242 19732 31260
rect 19224 31096 19234 31242
rect 19370 31096 19732 31242
rect 19224 31080 19732 31096
rect 18018 28354 18218 30744
rect 18018 28226 18024 28354
rect 18208 28226 18218 28354
rect 18018 28216 18218 28226
rect 15892 28141 16492 28200
rect 15892 28140 16493 28141
rect 15892 27900 16252 28140
rect 16492 27900 16493 28140
rect 15892 27899 16493 27900
rect 6672 25680 9952 27840
rect 15892 27661 16492 27899
rect 15892 27660 16493 27661
rect 15892 27420 16252 27660
rect 16492 27420 16493 27660
rect 15892 27419 16493 27420
rect 15892 27181 16492 27419
rect 15892 27180 16493 27181
rect 15892 26940 16252 27180
rect 16492 26940 16493 27180
rect 15892 26939 16493 26940
rect 15892 26880 16492 26939
rect 6672 1140 6972 25680
rect 6672 1020 6772 1140
rect 6892 1020 6972 1140
rect 6672 1000 6972 1020
rect 25312 1000 25612 43259
rect 28154 2392 28426 2408
rect 28154 2246 28342 2392
rect 28410 2246 28426 2392
rect 28154 2228 28426 2246
rect 28154 780 28334 2228
rect 27234 600 28334 780
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C1
timestamp 1711870259
transform 1 0 22222 0 1 40500
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C2
timestamp 1711870259
transform 1 0 22202 0 1 35060
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_LWYDVW  C3
timestamp 1711870259
transform 1 0 22202 0 1 29600
box -2650 -2600 2649 2600
use sky130_fd_pr__cap_mim_m3_1_WMZ6NR  C4
timestamp 1711870259
transform 1 0 12862 0 1 26540
box -3150 -2600 3149 2600
use high_voltage_logo  high_voltage_logo_0
timestamp 1711967973
transform 0 -1 6040 1 0 1262
box 0 0 42336 5768
use sky130_fd_pr__pfet_g5v0d10v5_AABD7U  M1
timestamp 1725649402
transform 1 0 28074 0 1 44395
box -308 -447 308 447
use sky130_fd_pr__pfet_g5v0d10v5_AABD7U  M2
timestamp 1725649402
transform 1 0 28074 0 1 43567
box -308 -447 308 447
use sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ  M3
timestamp 1725649402
transform -1 0 27438 0 1 44456
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ  M4
timestamp 1725649402
transform 1 0 27438 0 1 43628
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_RSSSV2  M8
timestamp 1717238374
transform 1 0 24330 0 1 3949
box -4258 -339 4258 339
use sky130_fd_pr__pfet_g5v0d10v5_RSSSV2  M9
timestamp 1717238374
transform 1 0 24330 0 1 2835
box -4258 -339 4258 339
use sky130_fd_pr__pfet_g5v0d10v5_RSSSV2  M10
timestamp 1717238374
transform 1 0 24330 0 1 1739
box -4258 -339 4258 339
use sky130_fd_pr__diode_pd2nw_11v0_AZAYX8  sky130_fd_pr__diode_pd2nw_11v0_AZAYX8_1
timestamp 1725619700
transform 1 0 18530 0 1 42186
box -478 -478 478 478
use sky130_fd_pr__diode_pd2nw_11v0_AZAYX8  sky130_fd_pr__diode_pd2nw_11v0_AZAYX8_2
timestamp 1725619700
transform 1 0 18538 0 1 36564
box -478 -478 478 478
use sky130_fd_pr__diode_pd2nw_11v0_AZAYX8  sky130_fd_pr__diode_pd2nw_11v0_AZAYX8_3
timestamp 1725619700
transform 1 0 18532 0 1 31156
box -478 -478 478 478
use sky130_fd_pr__diode_pd2nw_11v0_AZAYX8  sky130_fd_pr__diode_pd2nw_11v0_AZAYX8_4
timestamp 1725619700
transform 1 0 18532 0 1 27872
box -478 -478 478 478
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 25312 1000 25612 44152 1 FreeSans 2 0 0 0 VAPWR
port 51 nsew power bidirectional
flabel metal4 6672 1000 6972 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 6072 1000 6372 44152 1 FreeSans 2 0 0 0 VDPWR
port 53 nsew power bidirectional
flabel metal1 27632 43980 27692 44100 0 FreeSans 320 90 0 0 clka
flabel metal1 27552 42960 27612 43560 0 FreeSans 320 90 0 0 clkb
flabel metal2 19192 37800 19372 42120 0 FreeSans 1600 0 0 0 stage1
flabel metal2 19192 32400 19372 36480 0 FreeSans 1600 0 0 0 stage2
flabel metal3 16252 21660 16492 23880 0 FreeSans 1600 0 0 0 vout
flabel metal2 19208 28800 19388 31080 0 FreeSans 1600 0 0 0 stage3
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
