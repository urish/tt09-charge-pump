* NGSPICE file created from tt_um_urish_charge_pump.ext - technology: sky130A

.subckt tt_um_urish_charge_pump clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VPWR VGND
X0 clka clk.t0 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.45
X1 stage2.t4 clkb.t0 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X2 ua[0].t3 VGND.t3 VGND.t4 ua[0].t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=40
X3 stage3.t3 stage2.t1 stage2.t3 stage2.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=8
X4 VGND.t5 vout sky130_fd_pr__cap_mim_m3_1 l=25 w=30
X5 stage3.t4 clka.t0 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X6 clkb.t2 clka VGND.t2 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.45
X7 VPWR.t1 clk.t1 clka VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.45
X8 ua[0].t1 ua[0].t0 vout.t1 vout.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=40
X9 stage3.t2 stage3.t0 vout stage3.t1 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=8
X10 stage2.t0 stage1.t0 stage1.t2 stage1.t1 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=8
X11 stage1.t3 VPWR.t2 VPWR.t4 VPWR.t3 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=2.03 ps=14.58 w=7 l=8
X12 stage1.t4 clka.t1 sky130_fd_pr__cap_mim_m3_1 l=25 w=25
X13 VPWR.t5 clka.t2 clkb.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.45
R0 clk.n0 clk.t1 276.433
R1 clk.n0 clk.t0 244.831
R2 clk.n1 clk.n0 16.3372
R3 clk clk.n1 0.0952833
R4 clk.n1 clk 0.0189314
R5 VGND.n13 VGND.n9 2479.88
R6 VGND.n13 VGND.n10 2479.88
R7 VGND.n25 VGND.n9 2479.88
R8 VGND.n25 VGND.n10 2479.88
R9 VGND.n24 VGND.n18 2479.88
R10 VGND.n18 VGND.n14 2479.88
R11 VGND.n16 VGND.n14 2479.88
R12 VGND.n24 VGND.n16 2479.88
R13 VGND.n49 VGND.t4 660.787
R14 VGND.n15 VGND.n11 404.274
R15 VGND.n17 VGND.n11 404.274
R16 VGND.n26 VGND.n25 195
R17 VGND.n25 VGND.t0 195
R18 VGND.n13 VGND.n12 195
R19 VGND.t0 VGND.n13 195
R20 VGND.n24 VGND.n23 195
R21 VGND.t0 VGND.n24 195
R22 VGND.n20 VGND.n14 195
R23 VGND.t0 VGND.n14 195
R24 VGND.n12 VGND.n8 161.13
R25 VGND.n12 VGND.n7 161.13
R26 VGND.n26 VGND.n8 161.13
R27 VGND.n23 VGND.n19 161.13
R28 VGND.n20 VGND.n19 161.13
R29 VGND.n21 VGND.n20 161.13
R30 VGND.n27 VGND.n26 153.601
R31 VGND.n23 VGND.n22 139.294
R32 VGND.n10 VGND.n7 117.001
R33 VGND.n17 VGND.n10 117.001
R34 VGND.n9 VGND.n8 117.001
R35 VGND.n15 VGND.n9 117.001
R36 VGND.n19 VGND.n16 117.001
R37 VGND.n16 VGND.n15 117.001
R38 VGND.n21 VGND.n18 117.001
R39 VGND.n18 VGND.n17 117.001
R40 VGND.n6 VGND.t2 84.0308
R41 VGND.n28 VGND.t1 83.9547
R42 VGND.n50 VGND.n49 26.0302
R43 VGND.n22 VGND.n21 21.8358
R44 VGND.n28 VGND.n27 9.3005
R45 VGND.n22 VGND.n6 9.3005
R46 VGND.n27 VGND.n7 7.52991
R47 VGND.n49 VGND.t3 7.28674
R48 VGND.t0 VGND.n11 5.7035
R49 VGND.n29 VGND.n6 5.60682
R50 VGND.n29 VGND.n28 5.50342
R51 VGND.n47 VGND 4.20543
R52 VGND.n51 VGND.n50 3.8545
R53 VGND.n30 VGND.n29 3.05557
R54 VGND.n47 VGND.n46 2.62623
R55 VGND VGND.n51 0.365382
R56 VGND.n0 uio_oe[7] 0.32762
R57 VGND.n46 uio_oe[0] 0.213567
R58 VGND.n30 uo_out[0] 0.1979
R59 VGND.n31 uo_out[1] 0.1979
R60 VGND.n32 uo_out[2] 0.1979
R61 VGND.n33 uo_out[3] 0.1979
R62 VGND.n34 uo_out[4] 0.1979
R63 VGND.n35 uo_out[5] 0.1979
R64 VGND.n36 uo_out[6] 0.1979
R65 VGND.n37 uo_out[7] 0.1979
R66 VGND.n38 uio_out[0] 0.1979
R67 VGND.n39 uio_out[1] 0.1979
R68 VGND.n40 uio_out[2] 0.1979
R69 VGND.n41 uio_out[3] 0.1979
R70 VGND.n42 uio_out[4] 0.1979
R71 VGND.n43 uio_out[5] 0.1979
R72 VGND.n44 uio_out[6] 0.1979
R73 VGND.n45 uio_out[7] 0.1979
R74 VGND.n5 uio_oe[1] 0.1979
R75 VGND.n4 uio_oe[2] 0.1979
R76 VGND.n3 uio_oe[3] 0.1979
R77 VGND.n2 uio_oe[4] 0.1979
R78 VGND.n1 uio_oe[5] 0.1979
R79 VGND.n0 uio_oe[6] 0.1979
R80 VGND.n5 VGND.n4 0.13022
R81 VGND.n4 VGND.n3 0.13022
R82 VGND.n3 VGND.n2 0.13022
R83 VGND.n2 VGND.n1 0.13022
R84 VGND.n1 VGND.n0 0.13022
R85 VGND.n31 VGND.n30 0.13022
R86 VGND.n32 VGND.n31 0.13022
R87 VGND.n33 VGND.n32 0.13022
R88 VGND.n34 VGND.n33 0.13022
R89 VGND.n35 VGND.n34 0.13022
R90 VGND.n36 VGND.n35 0.13022
R91 VGND.n37 VGND.n36 0.13022
R92 VGND.n38 VGND.n37 0.13022
R93 VGND.n39 VGND.n38 0.13022
R94 VGND.n40 VGND.n39 0.13022
R95 VGND.n41 VGND.n40 0.13022
R96 VGND.n42 VGND.n41 0.13022
R97 VGND.n43 VGND.n42 0.13022
R98 VGND.n44 VGND.n43 0.13022
R99 VGND.n45 VGND.n44 0.13022
R100 VGND.n46 VGND.n45 0.1133
R101 VGND.n46 VGND.n5 0.07664
R102 VGND.n48 VGND.t5 0.0297714
R103 VGND.n48 VGND.n47 0.0164673
R104 VGND.n51 VGND.n48 0.0164673
R105 VGND.n50 VGND 0.0130333
R106 clka clka.t2 276.433
R107 clka.n0 clka.t0 19.2376
R108 clka.n0 clka.t1 10.2333
R109 clka clka.n0 6.03696
R110 stage2.n7 stage2.n2 10330.9
R111 stage2.n6 stage2.n5 10330.9
R112 stage2.n5 stage2.t2 1841.91
R113 stage2.n7 stage2.n3 1841.91
R114 stage2.n8 stage2.n1 671.247
R115 stage2.n4 stage2.n1 671.247
R116 stage2.n4 stage2.n0 671.247
R117 stage2.t3 stage2.n8 360.659
R118 stage2.t3 stage2.n0 281.224
R119 stage2.t3 stage2.t1 31.6676
R120 stage2.n8 stage2.n7 25.4353
R121 stage2.n5 stage2.n4 25.4353
R122 stage2.n6 stage2.n1 23.4005
R123 stage2.n2 stage2.n0 23.4005
R124 stage2.t2 stage2.n2 19.1855
R125 stage2.n3 stage2.n6 19.1855
R126 stage2.t4 stage2.t0 13.1042
R127 stage2.n3 stage2.t2 8.34551
R128 stage2.t3 stage2.t4 8.27133
R129 clkb clkb.t1 167.643
R130 clkb clkb.t2 83.7335
R131 clkb clkb.t0 9.32862
R132 ua[0].n11 ua[0].n10 8605.04
R133 ua[0].n8 ua[0].n5 8605.04
R134 ua[0].n5 ua[0].n4 3489.23
R135 ua[0].n10 ua[0].n9 3489.23
R136 ua[0].n12 ua[0].n3 1652.71
R137 ua[0].n7 ua[0].n3 1652.71
R138 ua[0].n13 ua[0].n12 1525.46
R139 ua[0].n7 ua[0].n6 1525.46
R140 ua[0].n0 ua[0].t1 660.448
R141 ua[0].n1 ua[0].t3 660.24
R142 ua[0].n13 ua[0].n2 127.248
R143 ua[0].n6 ua[0].n2 127.248
R144 ua[0].n5 ua[0].n2 37.0005
R145 ua[0].n10 ua[0].n3 37.0005
R146 ua[0].n0 ua[0].t0 13.0329
R147 ua[0].n6 ua[0].n1 9.98434
R148 ua[0].n14 ua[0].n13 9.3005
R149 ua[0] ua[0].n15 6.46994
R150 ua[0].n12 ua[0].n11 1.54217
R151 ua[0].n8 ua[0].n7 1.54217
R152 ua[0].n15 ua[0].n0 1.08544
R153 ua[0].n11 ua[0].n4 0.917376
R154 ua[0].n9 ua[0].n8 0.917376
R155 ua[0].n15 ua[0].n14 0.899115
R156 ua[0].n14 ua[0].n1 0.684342
R157 ua[0].n9 ua[0].t2 0.626126
R158 ua[0].t2 ua[0].n4 0.626126
R159 stage3.n8 stage3.n3 10330.9
R160 stage3.n7 stage3.n4 10330.9
R161 stage3.n19 stage3.n18 6978.85
R162 stage3.n18 stage3.n17 6978.85
R163 stage3.n17 stage3.n14 6978.85
R164 stage3.n19 stage3.n14 6978.85
R165 stage3.n20 stage3.n13 3802.7
R166 stage3.n16 stage3.n13 3802.7
R167 stage3.n16 stage3.n12 3802.7
R168 stage3.n20 stage3.n12 3802.7
R169 stage3.t1 stage3.n3 1841.91
R170 stage3.n5 stage3.n4 1841.91
R171 stage3.n21 stage3.n11 890.354
R172 stage3.n15 stage3.n11 890.354
R173 stage3.n15 stage3.n10 890.354
R174 stage3.n9 stage3.n2 671.247
R175 stage3.n6 stage3.n2 671.247
R176 stage3.n6 stage3.n1 671.247
R177 stage3.t4 stage3.n10 549.836
R178 stage3.n0 stage3.n1 358.776
R179 stage3.n0 stage3.n9 292.894
R180 stage3.t4 stage3.n21 291.954
R181 stage3.t4 stage3.t0 31.798
R182 stage3.n3 stage3.n2 25.4353
R183 stage3.n4 stage3.n1 25.4353
R184 stage3.n9 stage3.n8 23.4005
R185 stage3.n7 stage3.n6 23.4005
R186 stage3.n8 stage3.n5 19.1855
R187 stage3.t1 stage3.n7 19.1855
R188 stage3.t4 stage3.t2 13.8222
R189 stage3.t4 stage3.t3 13.743
R190 stage3.t4 stage3.n0 9.00675
R191 stage3.n5 stage3.t1 8.34551
R192 stage3.n13 stage3.n11 5.78175
R193 stage3.n18 stage3.n13 5.78175
R194 stage3.n12 stage3.n10 5.78175
R195 stage3.n14 stage3.n12 5.78175
R196 stage3.n21 stage3.n20 5.28621
R197 stage3.n20 stage3.n19 5.28621
R198 stage3.n16 stage3.n15 5.28621
R199 stage3.n17 stage3.n16 5.28621
R200 vout.n0 vout.t1 660.668
R201 vout vout.n0 12.7263
R202 vout.n0 vout.t0 640.452
R203 VPWR.n32 VPWR.n26 10330.9
R204 VPWR.n30 VPWR.n29 10330.9
R205 VPWR.n43 VPWR.n40 6978.85
R206 VPWR.n45 VPWR.n40 6978.85
R207 VPWR.n44 VPWR.n43 6978.85
R208 VPWR.n45 VPWR.n44 6978.85
R209 VPWR.n42 VPWR.n38 3802.7
R210 VPWR.n46 VPWR.n38 3802.7
R211 VPWR.n42 VPWR.n39 3802.7
R212 VPWR.n46 VPWR.n39 3802.7
R213 VPWR.n29 VPWR.n28 1841.91
R214 VPWR.n32 VPWR.n31 1841.91
R215 VPWR.n16 VPWR.n5 1718.82
R216 VPWR.n12 VPWR.n5 1718.82
R217 VPWR.n16 VPWR.n6 1718.82
R218 VPWR.n12 VPWR.n6 1718.82
R219 VPWR.n10 VPWR.n3 1718.82
R220 VPWR.n10 VPWR.n4 1718.82
R221 VPWR.n18 VPWR.n4 1718.82
R222 VPWR.n18 VPWR.n3 1718.82
R223 VPWR.n47 VPWR.n37 890.354
R224 VPWR.n41 VPWR.n37 890.354
R225 VPWR.n41 VPWR.n36 890.354
R226 VPWR.n33 VPWR.n25 671.247
R227 VPWR.n27 VPWR.n25 671.247
R228 VPWR.n27 VPWR.n24 671.247
R229 VPWR.n48 VPWR.n47 539.282
R230 VPWR.n34 VPWR.n33 354.26
R231 VPWR.n48 VPWR.n36 303.988
R232 VPWR.n34 VPWR.n24 297.413
R233 VPWR.n13 VPWR.n8 183.341
R234 VPWR.n15 VPWR.n14 183.341
R235 VPWR.n14 VPWR.n13 183.341
R236 VPWR.n9 VPWR.n1 183.341
R237 VPWR.n9 VPWR.n2 183.341
R238 VPWR.n19 VPWR.n2 183.341
R239 VPWR.n20 VPWR.n1 169.036
R240 VPWR.n0 VPWR.t1 167.94
R241 VPWR.n21 VPWR.t5 167.881
R242 VPWR.n8 VPWR.n7 160.754
R243 VPWR.n17 VPWR.t0 121.004
R244 VPWR.n11 VPWR.t0 121.004
R245 VPWR.n14 VPWR.n6 61.6672
R246 VPWR.n6 VPWR.t0 61.6672
R247 VPWR.n8 VPWR.n5 61.6672
R248 VPWR.n5 VPWR.t0 61.6672
R249 VPWR.n3 VPWR.n1 61.6672
R250 VPWR.t0 VPWR.n3 61.6672
R251 VPWR.n4 VPWR.n2 61.6672
R252 VPWR.t0 VPWR.n4 61.6672
R253 VPWR.n23 VPWR.t2 31.8306
R254 VPWR.n13 VPWR.n12 26.4291
R255 VPWR.n12 VPWR.n11 26.4291
R256 VPWR.n16 VPWR.n15 26.4291
R257 VPWR.n17 VPWR.n16 26.4291
R258 VPWR.n10 VPWR.n9 26.4291
R259 VPWR.n11 VPWR.n10 26.4291
R260 VPWR.n19 VPWR.n18 26.4291
R261 VPWR.n18 VPWR.n17 26.4291
R262 VPWR.n33 VPWR.n32 25.4353
R263 VPWR.n29 VPWR.n27 25.4353
R264 VPWR.n30 VPWR.n25 23.4005
R265 VPWR.n26 VPWR.n24 23.4005
R266 VPWR.n15 VPWR.n7 22.5887
R267 VPWR.n28 VPWR.n26 19.1855
R268 VPWR.n31 VPWR.n30 19.1855
R269 VPWR.n20 VPWR.n19 14.3064
R270 VPWR.n23 VPWR.t4 13.9149
R271 VPWR.n7 VPWR.n0 9.3005
R272 VPWR.n21 VPWR.n20 9.3005
R273 VPWR VPWR.n50 7.20367
R274 VPWR.n50 VPWR.n22 7.05903
R275 VPWR.n47 VPWR.n46 5.78175
R276 VPWR.n46 VPWR.n45 5.78175
R277 VPWR.n42 VPWR.n41 5.78175
R278 VPWR.n43 VPWR.n42 5.78175
R279 VPWR.n39 VPWR.n37 5.28621
R280 VPWR.n44 VPWR.n39 5.28621
R281 VPWR.n38 VPWR.n36 5.28621
R282 VPWR.n40 VPWR.n38 5.28621
R283 VPWR.n35 VPWR.n34 4.6505
R284 VPWR.n31 VPWR.t3 4.17301
R285 VPWR.n28 VPWR.t3 4.17301
R286 VPWR.n50 VPWR.n49 3.42531
R287 VPWR.n49 VPWR.n48 3.1005
R288 VPWR.n22 VPWR.n0 1.46092
R289 VPWR.n49 VPWR.n35 0.15675
R290 VPWR.n35 VPWR.n23 0.0551875
R291 VPWR.n22 VPWR.n21 0.00258333
R292 stage1.n7 stage1.n2 10330.9
R293 stage1.n6 stage1.n5 10330.9
R294 stage1.n16 stage1.n13 6978.85
R295 stage1.n18 stage1.n13 6978.85
R296 stage1.n17 stage1.n16 6978.85
R297 stage1.n18 stage1.n17 6978.85
R298 stage1.n15 stage1.n11 3802.7
R299 stage1.n19 stage1.n11 3802.7
R300 stage1.n15 stage1.n12 3802.7
R301 stage1.n19 stage1.n12 3802.7
R302 stage1.n5 stage1.t1 1841.91
R303 stage1.n7 stage1.n3 1841.91
R304 stage1.n20 stage1.n10 890.354
R305 stage1.n14 stage1.n10 890.354
R306 stage1.n14 stage1.n9 890.354
R307 stage1.n8 stage1.n1 671.247
R308 stage1.n4 stage1.n1 671.247
R309 stage1.n4 stage1.n0 671.247
R310 stage1.t2 stage1.n20 572.424
R311 stage1.t2 stage1.n8 360.659
R312 stage1.t2 stage1.n0 281.224
R313 stage1.t2 stage1.n9 269.365
R314 stage1.t2 stage1.t0 31.6676
R315 stage1.n8 stage1.n7 25.4353
R316 stage1.n5 stage1.n4 25.4353
R317 stage1.n6 stage1.n1 23.4005
R318 stage1.n2 stage1.n0 23.4005
R319 stage1.t1 stage1.n2 19.1855
R320 stage1.n3 stage1.n6 19.1855
R321 stage1.t4 stage1.t3 13.5661
R322 stage1.t2 stage1.t4 9.94633
R323 stage1.n3 stage1.t1 8.34551
R324 stage1.n20 stage1.n19 5.78175
R325 stage1.n19 stage1.n18 5.78175
R326 stage1.n15 stage1.n14 5.78175
R327 stage1.n16 stage1.n15 5.78175
R328 stage1.n12 stage1.n10 5.28621
R329 stage1.n17 stage1.n12 5.28621
R330 stage1.n11 stage1.n9 5.28621
R331 stage1.n13 stage1.n11 5.28621
C0 clk ui_in[1] 2.07e-20
C1 uio_in[1] uio_in[2] 0.031023f
C2 clka VPWR 5.07751f
C3 clka dw_19800_30000# 0.101107f
C4 ui_in[5] ui_in[6] 0.031023f
C5 uio_in[5] uio_in[4] 0.031023f
C6 ui_in[6] VPWR 1.03e-19
C7 clkb VPWR 1.72951f
C8 uio_in[3] VPWR 1.03e-19
C9 uio_in[3] uio_in[2] 0.031023f
C10 clka clkb 2.835f
C11 m2_3592_35982# m2_2808_33406# 0.0711f
C12 ui_in[2] VPWR 1.03e-19
C13 ui_in[1] VPWR 1.03e-19
C14 m2_3592_35982# m2_3592_39062# 0.162853f
C15 m2_3592_15598# m2_2584_17838# 0.151985f
C16 rst_n clk 0.031944f
C17 ui_in[0] ui_in[1] 0.031023f
C18 m2_3648_12070# m2_2864_8934# 0.135204f
C19 ui_in[3] ui_in[4] 0.031023f
C20 ui_in[7] VPWR 1.03e-19
C21 ui_in[7] uio_in[0] 0.031023f
C22 m2_1800_4342# ua[6] 0.004395f
C23 ui_in[3] VPWR 1.03e-19
C24 uio_in[4] VPWR 1.03e-19
C25 uio_in[5] VPWR 1.03e-19
C26 uio_in[5] uio_in[6] 0.031023f
C27 m2_3592_39062# m2_3592_42086# 0.130452f
C28 ena clk 0.034743f
C29 m2_2584_29654# m2_2808_33406# 0.041637f
C30 clk VPWR 0.404729f
C31 m2_2472_13022# m2_2864_8934# 0.017782f
C32 m2_1800_4342# m2_3592_4230# 0.559432f
C33 ui_in[0] clk 9.82e-20
C34 clka clk 0.366934f
C35 ui_in[6] ui_in[7] 0.031023f
C36 rst_n VPWR 1.03e-19
C37 ui_in[2] ui_in[1] 0.031023f
C38 uio_in[6] uio_in[7] 0.031023f
C39 ui_in[0] rst_n 0.031023f
C40 vout ua[0] 12.5848f
C41 ui_in[5] ui_in[4] 0.031023f
C42 uio_in[3] uio_in[4] 0.031023f
C43 clka rst_n 3.03e-19
C44 m2_3592_15598# m2_3648_12070# 0.104769f
C45 vout VPWR 0.118949f
C46 ui_in[5] VPWR 1.03e-19
C47 m2_2472_13022# m2_3648_12070# 0.105624f
C48 ua[0] VPWR 0.268291f
C49 ua[0] ua[1] 0.001614f
C50 ui_in[4] VPWR 1.03e-19
C51 ui_in[2] ui_in[3] 0.031023f
C52 m2_2584_29654# m2_3592_27358# 0.091013f
C53 uio_in[1] VPWR 1.03e-19
C54 uio_in[0] VPWR 1.03e-19
C55 uio_in[1] uio_in[0] 0.031023f
C56 m2_1800_4342# m2_2864_8934# 0.00172f
C57 m2_2864_23326# m2_3592_27358# 0.138713f
C58 ui_in[0] VPWR 1.03e-19
C59 uio_in[2] VPWR 1.03e-19
C60 ua[1] VGND 0.145965f
C61 ua[2] VGND 0.148302f
C62 ua[3] VGND 0.148302f
C63 ua[4] VGND 0.148302f
C64 ua[5] VGND 0.148302f
C65 ua[6] VGND 0.142703f
C66 ua[7] VGND 0.146962f
C67 ena VGND 0.075936f
C68 rst_n VGND 0.04853f
C69 ui_in[0] VGND 0.048746f
C70 ui_in[1] VGND 0.048746f
C71 ui_in[2] VGND 0.048746f
C72 ui_in[3] VGND 0.048746f
C73 ui_in[4] VGND 0.048746f
C74 ui_in[5] VGND 0.048746f
C75 ui_in[6] VGND 0.048746f
C76 ui_in[7] VGND 0.048746f
C77 uio_in[0] VGND 0.048746f
C78 uio_in[1] VGND 0.048746f
C79 uio_in[2] VGND 0.048746f
C80 uio_in[3] VGND 0.048746f
C81 uio_in[4] VGND 0.048746f
C82 uio_in[5] VGND 0.048746f
C83 uio_in[6] VGND 0.048746f
C84 uio_in[7] VGND 0.079769f
C85 clk VGND 1.75558f
C86 ua[0] VGND 45.063232f
C87 VPWR VGND 49.884384f
C88 m2_3592_4230# VGND 2.41736f $ **FLOATING
C89 m2_1800_4342# VGND 11.662f $ **FLOATING
C90 m2_2864_8934# VGND 5.1283f $ **FLOATING
C91 m2_3648_12070# VGND 3.18023f $ **FLOATING
C92 m2_2472_13022# VGND 0.831538f $ **FLOATING
C93 m2_3592_15598# VGND 5.94344f $ **FLOATING
C94 m2_2584_17838# VGND 4.71527f $ **FLOATING
C95 m2_2864_23326# VGND 4.89346f $ **FLOATING
C96 m2_3592_27358# VGND 4.41841f $ **FLOATING
C97 m2_2584_29654# VGND 4.17312f $ **FLOATING
C98 m2_2808_33406# VGND 4.18017f $ **FLOATING
C99 m2_3592_35982# VGND 4.2612f $ **FLOATING
C100 m2_3592_39062# VGND 5.95916f $ **FLOATING
C101 m2_3592_42086# VGND 4.32567f $ **FLOATING
C102 clkb VGND 16.841198f
C103 clka VGND 32.061157f
C104 vout VGND 0.129604p
C105 dw_19800_30000# VGND 22.1302f $ **FLOATING
C106 stage1.t4 VGND 48.4045f
C107 stage1.t2 VGND 1.49534f
C108 stage1.t3 VGND 0.082135f
C109 stage1.t0 VGND 1.96445f
C110 stage1.n0 VGND 0.041838f
C111 stage1.n1 VGND 0.058955f
C112 stage1.n2 VGND 0.058955f
C113 stage1.t1 VGND 0.860174f
C114 stage1.n3 VGND 0.860174f
C115 stage1.n4 VGND 0.059019f
C116 stage1.n5 VGND 1.03182f
C117 stage1.n6 VGND 0.058955f
C118 stage1.n7 VGND 1.05319f
C119 stage1.n8 VGND 0.045369f
C120 stage1.n9 VGND 0.050911f
C121 stage1.n10 VGND 0.078034f
C122 stage1.n11 VGND 0.169751f
C123 stage1.n12 VGND 0.169751f
C124 stage1.n13 VGND 0.614204f
C125 stage1.n14 VGND 0.078084f
C126 stage1.n15 VGND 0.170037f
C127 stage1.n16 VGND 0.622947f
C128 stage1.n17 VGND 0.614204f
C129 stage1.n18 VGND 0.622947f
C130 stage1.n19 VGND 0.170037f
C131 stage1.n20 VGND 0.06418f
C132 VPWR.t1 VGND 0.003038f
C133 VPWR.n0 VGND 0.007327f
C134 VPWR.t5 VGND 0.003036f
C135 VPWR.n1 VGND 0.003132f
C136 VPWR.n2 VGND 0.003257f
C137 VPWR.n3 VGND 0.003257f
C138 VPWR.n4 VGND 0.003257f
C139 VPWR.t0 VGND 0.052347f
C140 VPWR.n5 VGND 0.003257f
C141 VPWR.n6 VGND 0.003257f
C142 VPWR.n7 VGND 0.00161f
C143 VPWR.n8 VGND 0.003059f
C144 VPWR.n9 VGND 0.003208f
C145 VPWR.n10 VGND 0.003208f
C146 VPWR.n11 VGND 0.040931f
C147 VPWR.n12 VGND 0.003208f
C148 VPWR.n13 VGND 0.003208f
C149 VPWR.n14 VGND 0.003257f
C150 VPWR.n15 VGND 0.001796f
C151 VPWR.n16 VGND 0.003208f
C152 VPWR.n17 VGND 0.040931f
C153 VPWR.n18 VGND 0.003208f
C154 VPWR.n19 VGND 0.001726f
C155 VPWR.n20 VGND 0.001607f
C156 VPWR.n21 VGND 0.004455f
C157 VPWR.n22 VGND 0.012893f
C158 VPWR.t2 VGND 0.385055f
C159 VPWR.t4 VGND 0.015767f
C160 VPWR.n23 VGND 0.140432f
C161 VPWR.n24 VGND 0.008313f
C162 VPWR.n25 VGND 0.011539f
C163 VPWR.n26 VGND 0.011539f
C164 VPWR.t3 VGND 0.33671f
C165 VPWR.n27 VGND 0.011551f
C166 VPWR.n29 VGND 0.201951f
C167 VPWR.n30 VGND 0.011539f
C168 VPWR.n32 VGND 0.206132f
C169 VPWR.n33 VGND 0.008813f
C170 VPWR.n34 VGND 0.006552f
C171 VPWR.n35 VGND 0.009005f
C172 VPWR.n36 VGND 0.01027f
C173 VPWR.n37 VGND 0.015273f
C174 VPWR.n38 VGND 0.033224f
C175 VPWR.n39 VGND 0.033224f
C176 VPWR.n40 VGND 0.120213f
C177 VPWR.n41 VGND 0.015283f
C178 VPWR.n42 VGND 0.03328f
C179 VPWR.n43 VGND 0.121925f
C180 VPWR.n44 VGND 0.120213f
C181 VPWR.n45 VGND 0.121925f
C182 VPWR.n46 VGND 0.03328f
C183 VPWR.n47 VGND 0.012283f
C184 VPWR.n48 VGND 0.009678f
C185 VPWR.n49 VGND 0.129525f
C186 VPWR.n50 VGND 1.41234f
C187 vout.t0 VGND 1.4301f
C188 vout.t1 VGND 0.00116f
C189 vout.n0 VGND 0.693297f
C190 stage3.n0 VGND 0.032636f
C191 stage3.t4 VGND 47.8291f
C192 stage3.t3 VGND 0.077522f
C193 stage3.t0 VGND 1.91766f
C194 stage3.t2 VGND 0.077969f
C195 stage3.n1 VGND 0.044103f
C196 stage3.n2 VGND 0.057545f
C197 stage3.n3 VGND 1.02688f
C198 stage3.n4 VGND 1.00606f
C199 stage3.t1 VGND 0.838692f
C200 stage3.n5 VGND 0.838692f
C201 stage3.n6 VGND 0.057482f
C202 stage3.n7 VGND 0.057482f
C203 stage3.n8 VGND 0.057482f
C204 stage3.n9 VGND 0.041221f
C205 stage3.n10 VGND 0.061605f
C206 stage3.n11 VGND 0.076134f
C207 stage3.n12 VGND 0.16579f
C208 stage3.n13 VGND 0.16579f
C209 stage3.n14 VGND 0.60739f
C210 stage3.n15 VGND 0.076085f
C211 stage3.n16 VGND 0.165511f
C212 stage3.n17 VGND 0.598865f
C213 stage3.n18 VGND 0.60739f
C214 stage3.n19 VGND 0.598865f
C215 stage3.n20 VGND 0.165511f
C216 stage3.n21 VGND 0.050586f
C217 ua[0].t1 VGND 0.005268f
C218 ua[0].t0 VGND 2.96209f
C219 ua[0].n0 VGND 0.263857f
C220 ua[0].t3 VGND 0.005265f
C221 ua[0].n1 VGND 0.025355f
C222 ua[0].n2 VGND 0.013735f
C223 ua[0].n3 VGND 0.173955f
C224 ua[0].n5 VGND 1.99399f
C225 ua[0].n6 VGND 0.087333f
C226 ua[0].n7 VGND 0.166073f
C227 ua[0].n8 VGND 0.293969f
C228 ua[0].t2 VGND 3.28704f
C229 ua[0].n10 VGND 1.99399f
C230 ua[0].n11 VGND 0.293969f
C231 ua[0].n12 VGND 0.166073f
C232 ua[0].n13 VGND 0.086792f
C233 ua[0].n14 VGND 0.014191f
C234 ua[0].n15 VGND 0.086114f
C235 clkb.t0 VGND 58.603302f
C236 clkb.t2 VGND 0.020864f
C237 clkb.t1 VGND 0.032902f
C238 stage2.t3 VGND 1.80979f
C239 stage2.t4 VGND 62.691597f
C240 stage2.t0 VGND 0.096294f
C241 stage2.t1 VGND 2.54782f
C242 stage2.n0 VGND 0.054262f
C243 stage2.n1 VGND 0.076462f
C244 stage2.n2 VGND 0.076462f
C245 stage2.t2 VGND 1.11561f
C246 stage2.n3 VGND 1.11561f
C247 stage2.n4 VGND 0.076546f
C248 stage2.n5 VGND 1.33824f
C249 stage2.n6 VGND 0.076462f
C250 stage2.n7 VGND 1.36594f
C251 stage2.n8 VGND 0.058842f
C252 clka.t2 VGND 0.080865f
C253 clka.t0 VGND 60.1965f
C254 clka.t1 VGND 58.862103f
C255 clka.n0 VGND 2.94109f
.ends

